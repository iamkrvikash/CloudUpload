VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_2_16_scn4m_subm
   CLASS BLOCK ;
   SIZE 206.7 BY 422.0 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  106.4 39.6 107.2 40.4 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  128.2 39.6 129.0 40.4 ;
      END
   END din0[1]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  62.8 350.6 63.6 351.4 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  62.8 372.6 63.6 373.4 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  62.8 390.6 63.6 391.4 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  62.8 412.6 63.6 413.4 ;
      END
   END addr0[3]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  7.6 8.6 8.4 9.4 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  7.6 30.6 8.4 31.4 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  51.7 9.5 52.3 10.1 ;
      END
   END clk0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER m2 ;
         RECT  185.1 109.8 185.9 112.8 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER m2 ;
         RECT  191.9 109.8 192.7 112.8 ;
      END
   END dout0[1]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER m3 ;
         RECT  173.9 360.0 174.7 360.8 ;
         LAYER m3 ;
         RECT  20.8 221.2 21.6 222.0 ;
         LAYER m3 ;
         RECT  195.1 71.2 195.9 72.0 ;
         LAYER m3 ;
         RECT  173.9 318.4 174.7 319.2 ;
         LAYER m3 ;
         RECT  7.6 182.0 8.4 182.8 ;
         LAYER m3 ;
         RECT  131.1 50.6 131.9 51.4 ;
         LAYER m3 ;
         RECT  75.2 99.6 76.0 100.4 ;
         LAYER m3 ;
         RECT  165.1 339.6 165.9 340.4 ;
         LAYER m3 ;
         RECT  201.1 235.2 201.9 236.0 ;
         LAYER m3 ;
         RECT  173.9 172.8 174.7 173.6 ;
         LAYER m3 ;
         RECT  201.1 276.8 201.9 277.6 ;
         LAYER m3 ;
         RECT  201.1 339.2 201.9 340.0 ;
         LAYER m3 ;
         RECT  189.9 122.6 190.7 123.4 ;
         LAYER m3 ;
         RECT  165.1 298.0 165.9 298.8 ;
         LAYER m3 ;
         RECT  7.6 221.2 8.4 222.0 ;
         LAYER m3 ;
         RECT  -0.4 19.6 0.4 20.4 ;
         LAYER m3 ;
         RECT  105.7 214.8 106.5 215.6 ;
         LAYER m3 ;
         RECT  173.9 193.6 174.7 194.4 ;
         LAYER m3 ;
         RECT  7.6 299.6 8.4 300.4 ;
         LAYER m3 ;
         RECT  149.6 339.6 150.4 340.4 ;
         LAYER m3 ;
         RECT  194.5 88.6 195.3 89.4 ;
         LAYER m3 ;
         RECT  165.1 235.6 165.9 236.4 ;
         LAYER m3 ;
         RECT  201.1 297.6 201.9 298.4 ;
         LAYER m3 ;
         RECT  173.9 235.2 174.7 236.0 ;
         LAYER m3 ;
         RECT  20.8 338.8 21.6 339.6 ;
         LAYER m3 ;
         RECT  188.3 71.2 189.1 72.0 ;
         LAYER m3 ;
         RECT  20.8 299.6 21.6 300.4 ;
         LAYER m3 ;
         RECT  196.7 122.6 197.5 123.4 ;
         LAYER m3 ;
         RECT  187.5 172.8 188.3 173.6 ;
         LAYER m3 ;
         RECT  173.9 297.6 174.7 298.4 ;
         LAYER m3 ;
         RECT  149.6 235.6 150.4 236.4 ;
         LAYER m3 ;
         RECT  105.7 277.2 106.5 278.0 ;
         LAYER m3 ;
         RECT  90.7 256.4 91.5 257.2 ;
         LAYER m3 ;
         RECT  75.2 139.6 76.0 140.4 ;
         LAYER m3 ;
         RECT  187.7 88.6 188.5 89.4 ;
         LAYER m3 ;
         RECT  201.1 193.6 201.9 194.4 ;
         LAYER m3 ;
         RECT  173.9 276.8 174.7 277.6 ;
         LAYER m3 ;
         RECT  187.5 360.0 188.3 360.8 ;
         LAYER m3 ;
         RECT  201.1 172.8 201.9 173.6 ;
         LAYER m3 ;
         RECT  173.9 256.0 174.7 256.8 ;
         LAYER m3 ;
         RECT  201.1 318.4 201.9 319.2 ;
         LAYER m3 ;
         RECT  188.0 156.8 188.8 157.6 ;
         LAYER m3 ;
         RECT  180.7 360.0 181.5 360.8 ;
         LAYER m3 ;
         RECT  165.1 318.8 165.9 319.6 ;
         LAYER m3 ;
         RECT  165.1 277.2 165.9 278.0 ;
         LAYER m3 ;
         RECT  194.8 156.8 195.6 157.6 ;
         LAYER m3 ;
         RECT  20.8 260.4 21.6 261.2 ;
         LAYER m3 ;
         RECT  75.2 19.6 76.0 20.4 ;
         LAYER m3 ;
         RECT  65.7 401.6 66.5 402.4 ;
         LAYER m3 ;
         RECT  173.9 214.4 174.7 215.2 ;
         LAYER m3 ;
         RECT  149.6 277.2 150.4 278.0 ;
         LAYER m3 ;
         RECT  165.1 194.0 165.9 194.8 ;
         LAYER m3 ;
         RECT  105.7 194.0 106.5 194.8 ;
         LAYER m3 ;
         RECT  149.6 214.8 150.4 215.6 ;
         LAYER m3 ;
         RECT  173.9 339.2 174.7 340.0 ;
         LAYER m3 ;
         RECT  90.7 277.2 91.5 278.0 ;
         LAYER m3 ;
         RECT  201.1 256.0 201.9 256.8 ;
         LAYER m3 ;
         RECT  180.7 172.8 181.5 173.6 ;
         LAYER m3 ;
         RECT  181.2 156.8 182.0 157.6 ;
         LAYER m3 ;
         RECT  7.6 260.4 8.4 261.2 ;
         LAYER m3 ;
         RECT  201.1 214.4 201.9 215.2 ;
         LAYER m3 ;
         RECT  20.8 182.0 21.6 182.8 ;
         LAYER m3 ;
         RECT  165.1 256.4 165.9 257.2 ;
         LAYER m3 ;
         RECT  65.7 361.6 66.5 362.4 ;
         LAYER m3 ;
         RECT  201.1 360.0 201.9 360.8 ;
         LAYER m3 ;
         RECT  109.3 50.6 110.1 51.4 ;
         LAYER m3 ;
         RECT  90.7 214.8 91.5 215.6 ;
         LAYER m3 ;
         RECT  194.3 172.8 195.1 173.6 ;
         LAYER m3 ;
         RECT  75.2 59.6 76.0 60.4 ;
         LAYER m3 ;
         RECT  149.6 256.4 150.4 257.2 ;
         LAYER m3 ;
         RECT  105.7 256.4 106.5 257.2 ;
         LAYER m3 ;
         RECT  90.7 194.0 91.5 194.8 ;
         LAYER m3 ;
         RECT  165.1 214.8 165.9 215.6 ;
         LAYER m3 ;
         RECT  7.6 338.8 8.4 339.6 ;
         LAYER m3 ;
         RECT  149.6 318.8 150.4 319.6 ;
         LAYER m3 ;
         RECT  194.3 360.0 195.1 360.8 ;
         LAYER m3 ;
         RECT  149.6 298.0 150.4 298.8 ;
         LAYER m3 ;
         RECT  149.6 194.0 150.4 194.8 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER m3 ;
         RECT  204.5 219.4 205.3 220.2 ;
         LAYER m3 ;
         RECT  204.5 251.0 205.3 251.8 ;
         LAYER m3 ;
         RECT  189.7 82.2 190.5 83.0 ;
         LAYER m3 ;
         RECT  20.8 280.0 21.6 280.8 ;
         LAYER m3 ;
         RECT  165.1 329.2 165.9 330.0 ;
         LAYER m3 ;
         RECT  149.6 266.8 150.4 267.6 ;
         LAYER m3 ;
         RECT  204.5 344.2 205.3 345.0 ;
         LAYER m3 ;
         RECT  195.1 77.8 195.9 78.6 ;
         LAYER m3 ;
         RECT  197.7 344.2 198.5 345.0 ;
         LAYER m3 ;
         RECT  177.3 261.0 178.1 261.8 ;
         LAYER m3 ;
         RECT  170.5 313.4 171.3 314.2 ;
         LAYER m3 ;
         RECT  177.3 251.0 178.1 251.8 ;
         LAYER m3 ;
         RECT  204.5 271.8 205.3 272.6 ;
         LAYER m3 ;
         RECT  170.5 281.8 171.3 282.6 ;
         LAYER m3 ;
         RECT  75.2 159.6 76.0 160.4 ;
         LAYER m3 ;
         RECT  149.6 246.0 150.4 246.8 ;
         LAYER m3 ;
         RECT  188.3 77.8 189.1 78.6 ;
         LAYER m3 ;
         RECT  170.5 271.8 171.3 272.6 ;
         LAYER m3 ;
         RECT  197.7 281.8 198.5 282.6 ;
         LAYER m3 ;
         RECT  165.1 308.4 165.9 309.2 ;
         LAYER m3 ;
         RECT  177.3 271.8 178.1 272.6 ;
         LAYER m3 ;
         RECT  165.1 246.0 165.9 246.8 ;
         LAYER m3 ;
         RECT  90.7 183.6 91.5 184.4 ;
         LAYER m3 ;
         RECT  197.7 167.8 198.5 168.6 ;
         LAYER m3 ;
         RECT  7.6 319.2 8.4 320.0 ;
         LAYER m3 ;
         RECT  204.5 281.8 205.3 282.6 ;
         LAYER m3 ;
         RECT  90.7 287.6 91.5 288.4 ;
         LAYER m3 ;
         RECT  165.1 183.6 165.9 184.4 ;
         LAYER m3 ;
         RECT  197.7 198.6 198.5 199.4 ;
         LAYER m3 ;
         RECT  177.3 230.2 178.1 231.0 ;
         LAYER m3 ;
         RECT  197.7 209.4 198.5 210.2 ;
         LAYER m3 ;
         RECT  90.7 225.2 91.5 226.0 ;
         LAYER m3 ;
         RECT  170.5 177.8 171.3 178.6 ;
         LAYER m3 ;
         RECT  184.1 167.8 184.9 168.6 ;
         LAYER m3 ;
         RECT  204.5 177.8 205.3 178.6 ;
         LAYER m3 ;
         RECT  105.7 204.4 106.5 205.2 ;
         LAYER m3 ;
         RECT  204.5 302.6 205.3 303.4 ;
         LAYER m3 ;
         RECT  197.7 188.6 198.5 189.4 ;
         LAYER m3 ;
         RECT  204.5 313.4 205.3 314.2 ;
         LAYER m3 ;
         RECT  177.3 219.4 178.1 220.2 ;
         LAYER m3 ;
         RECT  204.5 323.4 205.3 324.2 ;
         LAYER m3 ;
         RECT  170.5 334.2 171.3 335.0 ;
         LAYER m3 ;
         RECT  193.7 96.8 194.5 97.6 ;
         LAYER m3 ;
         RECT  170.5 219.4 171.3 220.2 ;
         LAYER m3 ;
         RECT  197.7 302.6 198.5 303.4 ;
         LAYER m3 ;
         RECT  197.7 219.4 198.5 220.2 ;
         LAYER m3 ;
         RECT  197.7 292.6 198.5 293.4 ;
         LAYER m3 ;
         RECT  186.9 96.8 187.7 97.6 ;
         LAYER m3 ;
         RECT  177.3 355.0 178.1 355.8 ;
         LAYER m3 ;
         RECT  197.7 323.4 198.5 324.2 ;
         LAYER m3 ;
         RECT  170.5 323.4 171.3 324.2 ;
         LAYER m3 ;
         RECT  204.5 209.4 205.3 210.2 ;
         LAYER m3 ;
         RECT  20.8 240.8 21.6 241.6 ;
         LAYER m3 ;
         RECT  177.3 209.4 178.1 210.2 ;
         LAYER m3 ;
         RECT  105.7 287.6 106.5 288.4 ;
         LAYER m3 ;
         RECT  165.1 225.2 165.9 226.0 ;
         LAYER m3 ;
         RECT  197.7 240.2 198.5 241.0 ;
         LAYER m3 ;
         RECT  7.6 201.6 8.4 202.4 ;
         LAYER m3 ;
         RECT  196.5 82.2 197.3 83.0 ;
         LAYER m3 ;
         RECT  170.5 261.0 171.3 261.8 ;
         LAYER m3 ;
         RECT  170.5 344.2 171.3 345.0 ;
         LAYER m3 ;
         RECT  65.7 421.6 66.5 422.4 ;
         LAYER m3 ;
         RECT  90.7 266.8 91.5 267.6 ;
         LAYER m3 ;
         RECT  190.9 167.8 191.7 168.6 ;
         LAYER m3 ;
         RECT  7.6 280.0 8.4 280.8 ;
         LAYER m3 ;
         RECT  204.5 355.0 205.3 355.8 ;
         LAYER m3 ;
         RECT  -0.4 39.6 0.4 40.4 ;
         LAYER m3 ;
         RECT  -0.4 -0.4 0.4 0.4 ;
         LAYER m3 ;
         RECT  177.3 292.6 178.1 293.4 ;
         LAYER m3 ;
         RECT  190.9 355.0 191.7 355.8 ;
         LAYER m3 ;
         RECT  177.3 323.4 178.1 324.2 ;
         LAYER m3 ;
         RECT  170.5 230.2 171.3 231.0 ;
         LAYER m3 ;
         RECT  170.5 302.6 171.3 303.4 ;
         LAYER m3 ;
         RECT  149.6 350.0 150.4 350.8 ;
         LAYER m3 ;
         RECT  105.7 266.8 106.5 267.6 ;
         LAYER m3 ;
         RECT  149.6 204.4 150.4 205.2 ;
         LAYER m3 ;
         RECT  149.6 308.4 150.4 309.2 ;
         LAYER m3 ;
         RECT  170.5 240.2 171.3 241.0 ;
         LAYER m3 ;
         RECT  197.7 251.0 198.5 251.8 ;
         LAYER m3 ;
         RECT  177.3 334.2 178.1 335.0 ;
         LAYER m3 ;
         RECT  177.3 198.6 178.1 199.4 ;
         LAYER m3 ;
         RECT  204.5 167.8 205.3 168.6 ;
         LAYER m3 ;
         RECT  184.1 355.0 184.9 355.8 ;
         LAYER m3 ;
         RECT  204.5 188.6 205.3 189.4 ;
         LAYER m3 ;
         RECT  131.1 30.6 131.9 31.4 ;
         LAYER m3 ;
         RECT  204.5 261.0 205.3 261.8 ;
         LAYER m3 ;
         RECT  20.8 319.2 21.6 320.0 ;
         LAYER m3 ;
         RECT  170.5 209.4 171.3 210.2 ;
         LAYER m3 ;
         RECT  7.6 162.4 8.4 163.2 ;
         LAYER m3 ;
         RECT  165.1 350.0 165.9 350.8 ;
         LAYER m3 ;
         RECT  170.5 251.0 171.3 251.8 ;
         LAYER m3 ;
         RECT  109.3 30.6 110.1 31.4 ;
         LAYER m3 ;
         RECT  197.7 230.2 198.5 231.0 ;
         LAYER m3 ;
         RECT  197.7 271.8 198.5 272.6 ;
         LAYER m3 ;
         RECT  177.3 281.8 178.1 282.6 ;
         LAYER m3 ;
         RECT  105.7 225.2 106.5 226.0 ;
         LAYER m3 ;
         RECT  170.5 355.0 171.3 355.8 ;
         LAYER m3 ;
         RECT  204.5 198.6 205.3 199.4 ;
         LAYER m3 ;
         RECT  177.3 167.8 178.1 168.6 ;
         LAYER m3 ;
         RECT  177.3 240.2 178.1 241.0 ;
         LAYER m3 ;
         RECT  105.7 183.6 106.5 184.4 ;
         LAYER m3 ;
         RECT  20.8 201.6 21.6 202.4 ;
         LAYER m3 ;
         RECT  170.5 188.6 171.3 189.4 ;
         LAYER m3 ;
         RECT  204.5 292.6 205.3 293.4 ;
         LAYER m3 ;
         RECT  190.9 136.0 191.7 136.8 ;
         LAYER m3 ;
         RECT  20.8 162.4 21.6 163.2 ;
         LAYER m3 ;
         RECT  65.7 381.6 66.5 382.4 ;
         LAYER m3 ;
         RECT  204.5 240.2 205.3 241.0 ;
         LAYER m3 ;
         RECT  177.3 313.4 178.1 314.2 ;
         LAYER m3 ;
         RECT  197.7 177.8 198.5 178.6 ;
         LAYER m3 ;
         RECT  7.6 240.8 8.4 241.6 ;
         LAYER m3 ;
         RECT  170.5 198.6 171.3 199.4 ;
         LAYER m3 ;
         RECT  165.1 287.6 165.9 288.4 ;
         LAYER m3 ;
         RECT  177.3 302.6 178.1 303.4 ;
         LAYER m3 ;
         RECT  165.1 266.8 165.9 267.6 ;
         LAYER m3 ;
         RECT  170.5 292.6 171.3 293.4 ;
         LAYER m3 ;
         RECT  197.7 334.2 198.5 335.0 ;
         LAYER m3 ;
         RECT  65.7 341.6 66.5 342.4 ;
         LAYER m3 ;
         RECT  165.1 204.4 165.9 205.2 ;
         LAYER m3 ;
         RECT  149.6 329.2 150.4 330.0 ;
         LAYER m3 ;
         RECT  177.3 344.2 178.1 345.0 ;
         LAYER m3 ;
         RECT  90.7 204.4 91.5 205.2 ;
         LAYER m3 ;
         RECT  75.2 119.6 76.0 120.4 ;
         LAYER m3 ;
         RECT  197.7 261.0 198.5 261.8 ;
         LAYER m3 ;
         RECT  149.6 225.2 150.4 226.0 ;
         LAYER m3 ;
         RECT  197.7 355.0 198.5 355.8 ;
         LAYER m3 ;
         RECT  177.3 177.8 178.1 178.6 ;
         LAYER m3 ;
         RECT  75.2 39.6 76.0 40.4 ;
         LAYER m3 ;
         RECT  197.7 136.0 198.5 136.8 ;
         LAYER m3 ;
         RECT  177.3 188.6 178.1 189.4 ;
         LAYER m3 ;
         RECT  149.6 183.6 150.4 184.4 ;
         LAYER m3 ;
         RECT  149.6 287.6 150.4 288.4 ;
         LAYER m3 ;
         RECT  204.5 230.2 205.3 231.0 ;
         LAYER m3 ;
         RECT  204.5 334.2 205.3 335.0 ;
         LAYER m3 ;
         RECT  75.2 79.6 76.0 80.4 ;
         LAYER m3 ;
         RECT  197.7 313.4 198.5 314.2 ;
         LAYER m3 ;
         RECT  90.7 246.0 91.5 246.8 ;
         LAYER m3 ;
         RECT  75.2 -0.4 76.0 0.4 ;
         LAYER m3 ;
         RECT  105.7 246.0 106.5 246.8 ;
         LAYER m3 ;
         RECT  170.5 167.8 171.3 168.6 ;
      END
   END gnd
   OBS
   LAYER  m1 ;
      RECT  184.1 193.6 191.7 194.4 ;
      RECT  186.7 190.6 188.3 191.4 ;
      RECT  189.1 189.6 189.9 192.0 ;
      RECT  190.9 187.2 191.7 191.4 ;
      RECT  184.1 185.8 191.7 186.6 ;
      RECT  187.9 186.6 188.7 186.8 ;
      RECT  186.7 191.4 187.5 192.0 ;
      RECT  188.9 192.0 189.9 192.8 ;
      RECT  186.5 187.6 187.5 188.4 ;
      RECT  190.9 192.0 191.7 193.6 ;
      RECT  184.1 192.0 184.9 193.6 ;
      RECT  188.7 188.8 189.9 189.6 ;
      RECT  189.1 188.4 189.9 188.8 ;
      RECT  189.1 187.6 190.1 188.4 ;
      RECT  185.7 184.4 187.3 185.2 ;
      RECT  188.5 184.4 190.1 185.2 ;
      RECT  186.7 192.0 187.7 192.8 ;
      RECT  184.1 187.2 184.9 191.4 ;
      RECT  186.7 188.4 187.5 190.6 ;
      RECT  184.1 194.4 191.7 193.6 ;
      RECT  186.7 197.4 188.3 196.6 ;
      RECT  189.1 198.4 189.9 196.0 ;
      RECT  190.9 200.8 191.7 196.6 ;
      RECT  184.1 202.2 191.7 201.4 ;
      RECT  187.9 201.4 188.7 201.2 ;
      RECT  186.7 196.6 187.5 196.0 ;
      RECT  188.9 196.0 189.9 195.2 ;
      RECT  186.5 200.4 187.5 199.6 ;
      RECT  190.9 196.0 191.7 194.4 ;
      RECT  184.1 196.0 184.9 194.4 ;
      RECT  188.7 199.2 189.9 198.4 ;
      RECT  189.1 199.6 189.9 199.2 ;
      RECT  189.1 200.4 190.1 199.6 ;
      RECT  185.7 203.6 187.3 202.8 ;
      RECT  188.5 203.6 190.1 202.8 ;
      RECT  186.7 196.0 187.7 195.2 ;
      RECT  184.1 200.8 184.9 196.6 ;
      RECT  186.7 199.6 187.5 197.4 ;
      RECT  184.1 214.4 191.7 215.2 ;
      RECT  186.7 211.4 188.3 212.2 ;
      RECT  189.1 210.4 189.9 212.8 ;
      RECT  190.9 208.0 191.7 212.2 ;
      RECT  184.1 206.6 191.7 207.4 ;
      RECT  187.9 207.4 188.7 207.6 ;
      RECT  186.7 212.2 187.5 212.8 ;
      RECT  188.9 212.8 189.9 213.6 ;
      RECT  186.5 208.4 187.5 209.2 ;
      RECT  190.9 212.8 191.7 214.4 ;
      RECT  184.1 212.8 184.9 214.4 ;
      RECT  188.7 209.6 189.9 210.4 ;
      RECT  189.1 209.2 189.9 209.6 ;
      RECT  189.1 208.4 190.1 209.2 ;
      RECT  185.7 205.2 187.3 206.0 ;
      RECT  188.5 205.2 190.1 206.0 ;
      RECT  186.7 212.8 187.7 213.6 ;
      RECT  184.1 208.0 184.9 212.2 ;
      RECT  186.7 209.2 187.5 211.4 ;
      RECT  184.1 215.2 191.7 214.4 ;
      RECT  186.7 218.2 188.3 217.4 ;
      RECT  189.1 219.2 189.9 216.8 ;
      RECT  190.9 221.6 191.7 217.4 ;
      RECT  184.1 223.0 191.7 222.2 ;
      RECT  187.9 222.2 188.7 222.0 ;
      RECT  186.7 217.4 187.5 216.8 ;
      RECT  188.9 216.8 189.9 216.0 ;
      RECT  186.5 221.2 187.5 220.4 ;
      RECT  190.9 216.8 191.7 215.2 ;
      RECT  184.1 216.8 184.9 215.2 ;
      RECT  188.7 220.0 189.9 219.2 ;
      RECT  189.1 220.4 189.9 220.0 ;
      RECT  189.1 221.2 190.1 220.4 ;
      RECT  185.7 224.4 187.3 223.6 ;
      RECT  188.5 224.4 190.1 223.6 ;
      RECT  186.7 216.8 187.7 216.0 ;
      RECT  184.1 221.6 184.9 217.4 ;
      RECT  186.7 220.4 187.5 218.2 ;
      RECT  184.1 235.2 191.7 236.0 ;
      RECT  186.7 232.2 188.3 233.0 ;
      RECT  189.1 231.2 189.9 233.6 ;
      RECT  190.9 228.8 191.7 233.0 ;
      RECT  184.1 227.4 191.7 228.2 ;
      RECT  187.9 228.2 188.7 228.4 ;
      RECT  186.7 233.0 187.5 233.6 ;
      RECT  188.9 233.6 189.9 234.4 ;
      RECT  186.5 229.2 187.5 230.0 ;
      RECT  190.9 233.6 191.7 235.2 ;
      RECT  184.1 233.6 184.9 235.2 ;
      RECT  188.7 230.4 189.9 231.2 ;
      RECT  189.1 230.0 189.9 230.4 ;
      RECT  189.1 229.2 190.1 230.0 ;
      RECT  185.7 226.0 187.3 226.8 ;
      RECT  188.5 226.0 190.1 226.8 ;
      RECT  186.7 233.6 187.7 234.4 ;
      RECT  184.1 228.8 184.9 233.0 ;
      RECT  186.7 230.0 187.5 232.2 ;
      RECT  184.1 236.0 191.7 235.2 ;
      RECT  186.7 239.0 188.3 238.2 ;
      RECT  189.1 240.0 189.9 237.6 ;
      RECT  190.9 242.4 191.7 238.2 ;
      RECT  184.1 243.8 191.7 243.0 ;
      RECT  187.9 243.0 188.7 242.8 ;
      RECT  186.7 238.2 187.5 237.6 ;
      RECT  188.9 237.6 189.9 236.8 ;
      RECT  186.5 242.0 187.5 241.2 ;
      RECT  190.9 237.6 191.7 236.0 ;
      RECT  184.1 237.6 184.9 236.0 ;
      RECT  188.7 240.8 189.9 240.0 ;
      RECT  189.1 241.2 189.9 240.8 ;
      RECT  189.1 242.0 190.1 241.2 ;
      RECT  185.7 245.2 187.3 244.4 ;
      RECT  188.5 245.2 190.1 244.4 ;
      RECT  186.7 237.6 187.7 236.8 ;
      RECT  184.1 242.4 184.9 238.2 ;
      RECT  186.7 241.2 187.5 239.0 ;
      RECT  184.1 256.0 191.7 256.8 ;
      RECT  186.7 253.0 188.3 253.8 ;
      RECT  189.1 252.0 189.9 254.4 ;
      RECT  190.9 249.6 191.7 253.8 ;
      RECT  184.1 248.2 191.7 249.0 ;
      RECT  187.9 249.0 188.7 249.2 ;
      RECT  186.7 253.8 187.5 254.4 ;
      RECT  188.9 254.4 189.9 255.2 ;
      RECT  186.5 250.0 187.5 250.8 ;
      RECT  190.9 254.4 191.7 256.0 ;
      RECT  184.1 254.4 184.9 256.0 ;
      RECT  188.7 251.2 189.9 252.0 ;
      RECT  189.1 250.8 189.9 251.2 ;
      RECT  189.1 250.0 190.1 250.8 ;
      RECT  185.7 246.8 187.3 247.6 ;
      RECT  188.5 246.8 190.1 247.6 ;
      RECT  186.7 254.4 187.7 255.2 ;
      RECT  184.1 249.6 184.9 253.8 ;
      RECT  186.7 250.8 187.5 253.0 ;
      RECT  184.1 256.8 191.7 256.0 ;
      RECT  186.7 259.8 188.3 259.0 ;
      RECT  189.1 260.8 189.9 258.4 ;
      RECT  190.9 263.2 191.7 259.0 ;
      RECT  184.1 264.6 191.7 263.8 ;
      RECT  187.9 263.8 188.7 263.6 ;
      RECT  186.7 259.0 187.5 258.4 ;
      RECT  188.9 258.4 189.9 257.6 ;
      RECT  186.5 262.8 187.5 262.0 ;
      RECT  190.9 258.4 191.7 256.8 ;
      RECT  184.1 258.4 184.9 256.8 ;
      RECT  188.7 261.6 189.9 260.8 ;
      RECT  189.1 262.0 189.9 261.6 ;
      RECT  189.1 262.8 190.1 262.0 ;
      RECT  185.7 266.0 187.3 265.2 ;
      RECT  188.5 266.0 190.1 265.2 ;
      RECT  186.7 258.4 187.7 257.6 ;
      RECT  184.1 263.2 184.9 259.0 ;
      RECT  186.7 262.0 187.5 259.8 ;
      RECT  184.1 276.8 191.7 277.6 ;
      RECT  186.7 273.8 188.3 274.6 ;
      RECT  189.1 272.8 189.9 275.2 ;
      RECT  190.9 270.4 191.7 274.6 ;
      RECT  184.1 269.0 191.7 269.8 ;
      RECT  187.9 269.8 188.7 270.0 ;
      RECT  186.7 274.6 187.5 275.2 ;
      RECT  188.9 275.2 189.9 276.0 ;
      RECT  186.5 270.8 187.5 271.6 ;
      RECT  190.9 275.2 191.7 276.8 ;
      RECT  184.1 275.2 184.9 276.8 ;
      RECT  188.7 272.0 189.9 272.8 ;
      RECT  189.1 271.6 189.9 272.0 ;
      RECT  189.1 270.8 190.1 271.6 ;
      RECT  185.7 267.6 187.3 268.4 ;
      RECT  188.5 267.6 190.1 268.4 ;
      RECT  186.7 275.2 187.7 276.0 ;
      RECT  184.1 270.4 184.9 274.6 ;
      RECT  186.7 271.6 187.5 273.8 ;
      RECT  184.1 277.6 191.7 276.8 ;
      RECT  186.7 280.6 188.3 279.8 ;
      RECT  189.1 281.6 189.9 279.2 ;
      RECT  190.9 284.0 191.7 279.8 ;
      RECT  184.1 285.4 191.7 284.6 ;
      RECT  187.9 284.6 188.7 284.4 ;
      RECT  186.7 279.8 187.5 279.2 ;
      RECT  188.9 279.2 189.9 278.4 ;
      RECT  186.5 283.6 187.5 282.8 ;
      RECT  190.9 279.2 191.7 277.6 ;
      RECT  184.1 279.2 184.9 277.6 ;
      RECT  188.7 282.4 189.9 281.6 ;
      RECT  189.1 282.8 189.9 282.4 ;
      RECT  189.1 283.6 190.1 282.8 ;
      RECT  185.7 286.8 187.3 286.0 ;
      RECT  188.5 286.8 190.1 286.0 ;
      RECT  186.7 279.2 187.7 278.4 ;
      RECT  184.1 284.0 184.9 279.8 ;
      RECT  186.7 282.8 187.5 280.6 ;
      RECT  184.1 297.6 191.7 298.4 ;
      RECT  186.7 294.6 188.3 295.4 ;
      RECT  189.1 293.6 189.9 296.0 ;
      RECT  190.9 291.2 191.7 295.4 ;
      RECT  184.1 289.8 191.7 290.6 ;
      RECT  187.9 290.6 188.7 290.8 ;
      RECT  186.7 295.4 187.5 296.0 ;
      RECT  188.9 296.0 189.9 296.8 ;
      RECT  186.5 291.6 187.5 292.4 ;
      RECT  190.9 296.0 191.7 297.6 ;
      RECT  184.1 296.0 184.9 297.6 ;
      RECT  188.7 292.8 189.9 293.6 ;
      RECT  189.1 292.4 189.9 292.8 ;
      RECT  189.1 291.6 190.1 292.4 ;
      RECT  185.7 288.4 187.3 289.2 ;
      RECT  188.5 288.4 190.1 289.2 ;
      RECT  186.7 296.0 187.7 296.8 ;
      RECT  184.1 291.2 184.9 295.4 ;
      RECT  186.7 292.4 187.5 294.6 ;
      RECT  184.1 298.4 191.7 297.6 ;
      RECT  186.7 301.4 188.3 300.6 ;
      RECT  189.1 302.4 189.9 300.0 ;
      RECT  190.9 304.8 191.7 300.6 ;
      RECT  184.1 306.2 191.7 305.4 ;
      RECT  187.9 305.4 188.7 305.2 ;
      RECT  186.7 300.6 187.5 300.0 ;
      RECT  188.9 300.0 189.9 299.2 ;
      RECT  186.5 304.4 187.5 303.6 ;
      RECT  190.9 300.0 191.7 298.4 ;
      RECT  184.1 300.0 184.9 298.4 ;
      RECT  188.7 303.2 189.9 302.4 ;
      RECT  189.1 303.6 189.9 303.2 ;
      RECT  189.1 304.4 190.1 303.6 ;
      RECT  185.7 307.6 187.3 306.8 ;
      RECT  188.5 307.6 190.1 306.8 ;
      RECT  186.7 300.0 187.7 299.2 ;
      RECT  184.1 304.8 184.9 300.6 ;
      RECT  186.7 303.6 187.5 301.4 ;
      RECT  184.1 318.4 191.7 319.2 ;
      RECT  186.7 315.4 188.3 316.2 ;
      RECT  189.1 314.4 189.9 316.8 ;
      RECT  190.9 312.0 191.7 316.2 ;
      RECT  184.1 310.6 191.7 311.4 ;
      RECT  187.9 311.4 188.7 311.6 ;
      RECT  186.7 316.2 187.5 316.8 ;
      RECT  188.9 316.8 189.9 317.6 ;
      RECT  186.5 312.4 187.5 313.2 ;
      RECT  190.9 316.8 191.7 318.4 ;
      RECT  184.1 316.8 184.9 318.4 ;
      RECT  188.7 313.6 189.9 314.4 ;
      RECT  189.1 313.2 189.9 313.6 ;
      RECT  189.1 312.4 190.1 313.2 ;
      RECT  185.7 309.2 187.3 310.0 ;
      RECT  188.5 309.2 190.1 310.0 ;
      RECT  186.7 316.8 187.7 317.6 ;
      RECT  184.1 312.0 184.9 316.2 ;
      RECT  186.7 313.2 187.5 315.4 ;
      RECT  184.1 319.2 191.7 318.4 ;
      RECT  186.7 322.2 188.3 321.4 ;
      RECT  189.1 323.2 189.9 320.8 ;
      RECT  190.9 325.6 191.7 321.4 ;
      RECT  184.1 327.0 191.7 326.2 ;
      RECT  187.9 326.2 188.7 326.0 ;
      RECT  186.7 321.4 187.5 320.8 ;
      RECT  188.9 320.8 189.9 320.0 ;
      RECT  186.5 325.2 187.5 324.4 ;
      RECT  190.9 320.8 191.7 319.2 ;
      RECT  184.1 320.8 184.9 319.2 ;
      RECT  188.7 324.0 189.9 323.2 ;
      RECT  189.1 324.4 189.9 324.0 ;
      RECT  189.1 325.2 190.1 324.4 ;
      RECT  185.7 328.4 187.3 327.6 ;
      RECT  188.5 328.4 190.1 327.6 ;
      RECT  186.7 320.8 187.7 320.0 ;
      RECT  184.1 325.6 184.9 321.4 ;
      RECT  186.7 324.4 187.5 322.2 ;
      RECT  184.1 339.2 191.7 340.0 ;
      RECT  186.7 336.2 188.3 337.0 ;
      RECT  189.1 335.2 189.9 337.6 ;
      RECT  190.9 332.8 191.7 337.0 ;
      RECT  184.1 331.4 191.7 332.2 ;
      RECT  187.9 332.2 188.7 332.4 ;
      RECT  186.7 337.0 187.5 337.6 ;
      RECT  188.9 337.6 189.9 338.4 ;
      RECT  186.5 333.2 187.5 334.0 ;
      RECT  190.9 337.6 191.7 339.2 ;
      RECT  184.1 337.6 184.9 339.2 ;
      RECT  188.7 334.4 189.9 335.2 ;
      RECT  189.1 334.0 189.9 334.4 ;
      RECT  189.1 333.2 190.1 334.0 ;
      RECT  185.7 330.0 187.3 330.8 ;
      RECT  188.5 330.0 190.1 330.8 ;
      RECT  186.7 337.6 187.7 338.4 ;
      RECT  184.1 332.8 184.9 337.0 ;
      RECT  186.7 334.0 187.5 336.2 ;
      RECT  184.1 340.0 191.7 339.2 ;
      RECT  186.7 343.0 188.3 342.2 ;
      RECT  189.1 344.0 189.9 341.6 ;
      RECT  190.9 346.4 191.7 342.2 ;
      RECT  184.1 347.8 191.7 347.0 ;
      RECT  187.9 347.0 188.7 346.8 ;
      RECT  186.7 342.2 187.5 341.6 ;
      RECT  188.9 341.6 189.9 340.8 ;
      RECT  186.5 346.0 187.5 345.2 ;
      RECT  190.9 341.6 191.7 340.0 ;
      RECT  184.1 341.6 184.9 340.0 ;
      RECT  188.7 344.8 189.9 344.0 ;
      RECT  189.1 345.2 189.9 344.8 ;
      RECT  189.1 346.0 190.1 345.2 ;
      RECT  185.7 349.2 187.3 348.4 ;
      RECT  188.5 349.2 190.1 348.4 ;
      RECT  186.7 341.6 187.7 340.8 ;
      RECT  184.1 346.4 184.9 342.2 ;
      RECT  186.7 345.2 187.5 343.0 ;
      RECT  190.9 193.6 198.5 194.4 ;
      RECT  193.5 190.6 195.1 191.4 ;
      RECT  195.9 189.6 196.7 192.0 ;
      RECT  197.7 187.2 198.5 191.4 ;
      RECT  190.9 185.8 198.5 186.6 ;
      RECT  194.7 186.6 195.5 186.8 ;
      RECT  193.5 191.4 194.3 192.0 ;
      RECT  195.7 192.0 196.7 192.8 ;
      RECT  193.3 187.6 194.3 188.4 ;
      RECT  197.7 192.0 198.5 193.6 ;
      RECT  190.9 192.0 191.7 193.6 ;
      RECT  195.5 188.8 196.7 189.6 ;
      RECT  195.9 188.4 196.7 188.8 ;
      RECT  195.9 187.6 196.9 188.4 ;
      RECT  192.5 184.4 194.1 185.2 ;
      RECT  195.3 184.4 196.9 185.2 ;
      RECT  193.5 192.0 194.5 192.8 ;
      RECT  190.9 187.2 191.7 191.4 ;
      RECT  193.5 188.4 194.3 190.6 ;
      RECT  190.9 194.4 198.5 193.6 ;
      RECT  193.5 197.4 195.1 196.6 ;
      RECT  195.9 198.4 196.7 196.0 ;
      RECT  197.7 200.8 198.5 196.6 ;
      RECT  190.9 202.2 198.5 201.4 ;
      RECT  194.7 201.4 195.5 201.2 ;
      RECT  193.5 196.6 194.3 196.0 ;
      RECT  195.7 196.0 196.7 195.2 ;
      RECT  193.3 200.4 194.3 199.6 ;
      RECT  197.7 196.0 198.5 194.4 ;
      RECT  190.9 196.0 191.7 194.4 ;
      RECT  195.5 199.2 196.7 198.4 ;
      RECT  195.9 199.6 196.7 199.2 ;
      RECT  195.9 200.4 196.9 199.6 ;
      RECT  192.5 203.6 194.1 202.8 ;
      RECT  195.3 203.6 196.9 202.8 ;
      RECT  193.5 196.0 194.5 195.2 ;
      RECT  190.9 200.8 191.7 196.6 ;
      RECT  193.5 199.6 194.3 197.4 ;
      RECT  190.9 214.4 198.5 215.2 ;
      RECT  193.5 211.4 195.1 212.2 ;
      RECT  195.9 210.4 196.7 212.8 ;
      RECT  197.7 208.0 198.5 212.2 ;
      RECT  190.9 206.6 198.5 207.4 ;
      RECT  194.7 207.4 195.5 207.6 ;
      RECT  193.5 212.2 194.3 212.8 ;
      RECT  195.7 212.8 196.7 213.6 ;
      RECT  193.3 208.4 194.3 209.2 ;
      RECT  197.7 212.8 198.5 214.4 ;
      RECT  190.9 212.8 191.7 214.4 ;
      RECT  195.5 209.6 196.7 210.4 ;
      RECT  195.9 209.2 196.7 209.6 ;
      RECT  195.9 208.4 196.9 209.2 ;
      RECT  192.5 205.2 194.1 206.0 ;
      RECT  195.3 205.2 196.9 206.0 ;
      RECT  193.5 212.8 194.5 213.6 ;
      RECT  190.9 208.0 191.7 212.2 ;
      RECT  193.5 209.2 194.3 211.4 ;
      RECT  190.9 215.2 198.5 214.4 ;
      RECT  193.5 218.2 195.1 217.4 ;
      RECT  195.9 219.2 196.7 216.8 ;
      RECT  197.7 221.6 198.5 217.4 ;
      RECT  190.9 223.0 198.5 222.2 ;
      RECT  194.7 222.2 195.5 222.0 ;
      RECT  193.5 217.4 194.3 216.8 ;
      RECT  195.7 216.8 196.7 216.0 ;
      RECT  193.3 221.2 194.3 220.4 ;
      RECT  197.7 216.8 198.5 215.2 ;
      RECT  190.9 216.8 191.7 215.2 ;
      RECT  195.5 220.0 196.7 219.2 ;
      RECT  195.9 220.4 196.7 220.0 ;
      RECT  195.9 221.2 196.9 220.4 ;
      RECT  192.5 224.4 194.1 223.6 ;
      RECT  195.3 224.4 196.9 223.6 ;
      RECT  193.5 216.8 194.5 216.0 ;
      RECT  190.9 221.6 191.7 217.4 ;
      RECT  193.5 220.4 194.3 218.2 ;
      RECT  190.9 235.2 198.5 236.0 ;
      RECT  193.5 232.2 195.1 233.0 ;
      RECT  195.9 231.2 196.7 233.6 ;
      RECT  197.7 228.8 198.5 233.0 ;
      RECT  190.9 227.4 198.5 228.2 ;
      RECT  194.7 228.2 195.5 228.4 ;
      RECT  193.5 233.0 194.3 233.6 ;
      RECT  195.7 233.6 196.7 234.4 ;
      RECT  193.3 229.2 194.3 230.0 ;
      RECT  197.7 233.6 198.5 235.2 ;
      RECT  190.9 233.6 191.7 235.2 ;
      RECT  195.5 230.4 196.7 231.2 ;
      RECT  195.9 230.0 196.7 230.4 ;
      RECT  195.9 229.2 196.9 230.0 ;
      RECT  192.5 226.0 194.1 226.8 ;
      RECT  195.3 226.0 196.9 226.8 ;
      RECT  193.5 233.6 194.5 234.4 ;
      RECT  190.9 228.8 191.7 233.0 ;
      RECT  193.5 230.0 194.3 232.2 ;
      RECT  190.9 236.0 198.5 235.2 ;
      RECT  193.5 239.0 195.1 238.2 ;
      RECT  195.9 240.0 196.7 237.6 ;
      RECT  197.7 242.4 198.5 238.2 ;
      RECT  190.9 243.8 198.5 243.0 ;
      RECT  194.7 243.0 195.5 242.8 ;
      RECT  193.5 238.2 194.3 237.6 ;
      RECT  195.7 237.6 196.7 236.8 ;
      RECT  193.3 242.0 194.3 241.2 ;
      RECT  197.7 237.6 198.5 236.0 ;
      RECT  190.9 237.6 191.7 236.0 ;
      RECT  195.5 240.8 196.7 240.0 ;
      RECT  195.9 241.2 196.7 240.8 ;
      RECT  195.9 242.0 196.9 241.2 ;
      RECT  192.5 245.2 194.1 244.4 ;
      RECT  195.3 245.2 196.9 244.4 ;
      RECT  193.5 237.6 194.5 236.8 ;
      RECT  190.9 242.4 191.7 238.2 ;
      RECT  193.5 241.2 194.3 239.0 ;
      RECT  190.9 256.0 198.5 256.8 ;
      RECT  193.5 253.0 195.1 253.8 ;
      RECT  195.9 252.0 196.7 254.4 ;
      RECT  197.7 249.6 198.5 253.8 ;
      RECT  190.9 248.2 198.5 249.0 ;
      RECT  194.7 249.0 195.5 249.2 ;
      RECT  193.5 253.8 194.3 254.4 ;
      RECT  195.7 254.4 196.7 255.2 ;
      RECT  193.3 250.0 194.3 250.8 ;
      RECT  197.7 254.4 198.5 256.0 ;
      RECT  190.9 254.4 191.7 256.0 ;
      RECT  195.5 251.2 196.7 252.0 ;
      RECT  195.9 250.8 196.7 251.2 ;
      RECT  195.9 250.0 196.9 250.8 ;
      RECT  192.5 246.8 194.1 247.6 ;
      RECT  195.3 246.8 196.9 247.6 ;
      RECT  193.5 254.4 194.5 255.2 ;
      RECT  190.9 249.6 191.7 253.8 ;
      RECT  193.5 250.8 194.3 253.0 ;
      RECT  190.9 256.8 198.5 256.0 ;
      RECT  193.5 259.8 195.1 259.0 ;
      RECT  195.9 260.8 196.7 258.4 ;
      RECT  197.7 263.2 198.5 259.0 ;
      RECT  190.9 264.6 198.5 263.8 ;
      RECT  194.7 263.8 195.5 263.6 ;
      RECT  193.5 259.0 194.3 258.4 ;
      RECT  195.7 258.4 196.7 257.6 ;
      RECT  193.3 262.8 194.3 262.0 ;
      RECT  197.7 258.4 198.5 256.8 ;
      RECT  190.9 258.4 191.7 256.8 ;
      RECT  195.5 261.6 196.7 260.8 ;
      RECT  195.9 262.0 196.7 261.6 ;
      RECT  195.9 262.8 196.9 262.0 ;
      RECT  192.5 266.0 194.1 265.2 ;
      RECT  195.3 266.0 196.9 265.2 ;
      RECT  193.5 258.4 194.5 257.6 ;
      RECT  190.9 263.2 191.7 259.0 ;
      RECT  193.5 262.0 194.3 259.8 ;
      RECT  190.9 276.8 198.5 277.6 ;
      RECT  193.5 273.8 195.1 274.6 ;
      RECT  195.9 272.8 196.7 275.2 ;
      RECT  197.7 270.4 198.5 274.6 ;
      RECT  190.9 269.0 198.5 269.8 ;
      RECT  194.7 269.8 195.5 270.0 ;
      RECT  193.5 274.6 194.3 275.2 ;
      RECT  195.7 275.2 196.7 276.0 ;
      RECT  193.3 270.8 194.3 271.6 ;
      RECT  197.7 275.2 198.5 276.8 ;
      RECT  190.9 275.2 191.7 276.8 ;
      RECT  195.5 272.0 196.7 272.8 ;
      RECT  195.9 271.6 196.7 272.0 ;
      RECT  195.9 270.8 196.9 271.6 ;
      RECT  192.5 267.6 194.1 268.4 ;
      RECT  195.3 267.6 196.9 268.4 ;
      RECT  193.5 275.2 194.5 276.0 ;
      RECT  190.9 270.4 191.7 274.6 ;
      RECT  193.5 271.6 194.3 273.8 ;
      RECT  190.9 277.6 198.5 276.8 ;
      RECT  193.5 280.6 195.1 279.8 ;
      RECT  195.9 281.6 196.7 279.2 ;
      RECT  197.7 284.0 198.5 279.8 ;
      RECT  190.9 285.4 198.5 284.6 ;
      RECT  194.7 284.6 195.5 284.4 ;
      RECT  193.5 279.8 194.3 279.2 ;
      RECT  195.7 279.2 196.7 278.4 ;
      RECT  193.3 283.6 194.3 282.8 ;
      RECT  197.7 279.2 198.5 277.6 ;
      RECT  190.9 279.2 191.7 277.6 ;
      RECT  195.5 282.4 196.7 281.6 ;
      RECT  195.9 282.8 196.7 282.4 ;
      RECT  195.9 283.6 196.9 282.8 ;
      RECT  192.5 286.8 194.1 286.0 ;
      RECT  195.3 286.8 196.9 286.0 ;
      RECT  193.5 279.2 194.5 278.4 ;
      RECT  190.9 284.0 191.7 279.8 ;
      RECT  193.5 282.8 194.3 280.6 ;
      RECT  190.9 297.6 198.5 298.4 ;
      RECT  193.5 294.6 195.1 295.4 ;
      RECT  195.9 293.6 196.7 296.0 ;
      RECT  197.7 291.2 198.5 295.4 ;
      RECT  190.9 289.8 198.5 290.6 ;
      RECT  194.7 290.6 195.5 290.8 ;
      RECT  193.5 295.4 194.3 296.0 ;
      RECT  195.7 296.0 196.7 296.8 ;
      RECT  193.3 291.6 194.3 292.4 ;
      RECT  197.7 296.0 198.5 297.6 ;
      RECT  190.9 296.0 191.7 297.6 ;
      RECT  195.5 292.8 196.7 293.6 ;
      RECT  195.9 292.4 196.7 292.8 ;
      RECT  195.9 291.6 196.9 292.4 ;
      RECT  192.5 288.4 194.1 289.2 ;
      RECT  195.3 288.4 196.9 289.2 ;
      RECT  193.5 296.0 194.5 296.8 ;
      RECT  190.9 291.2 191.7 295.4 ;
      RECT  193.5 292.4 194.3 294.6 ;
      RECT  190.9 298.4 198.5 297.6 ;
      RECT  193.5 301.4 195.1 300.6 ;
      RECT  195.9 302.4 196.7 300.0 ;
      RECT  197.7 304.8 198.5 300.6 ;
      RECT  190.9 306.2 198.5 305.4 ;
      RECT  194.7 305.4 195.5 305.2 ;
      RECT  193.5 300.6 194.3 300.0 ;
      RECT  195.7 300.0 196.7 299.2 ;
      RECT  193.3 304.4 194.3 303.6 ;
      RECT  197.7 300.0 198.5 298.4 ;
      RECT  190.9 300.0 191.7 298.4 ;
      RECT  195.5 303.2 196.7 302.4 ;
      RECT  195.9 303.6 196.7 303.2 ;
      RECT  195.9 304.4 196.9 303.6 ;
      RECT  192.5 307.6 194.1 306.8 ;
      RECT  195.3 307.6 196.9 306.8 ;
      RECT  193.5 300.0 194.5 299.2 ;
      RECT  190.9 304.8 191.7 300.6 ;
      RECT  193.5 303.6 194.3 301.4 ;
      RECT  190.9 318.4 198.5 319.2 ;
      RECT  193.5 315.4 195.1 316.2 ;
      RECT  195.9 314.4 196.7 316.8 ;
      RECT  197.7 312.0 198.5 316.2 ;
      RECT  190.9 310.6 198.5 311.4 ;
      RECT  194.7 311.4 195.5 311.6 ;
      RECT  193.5 316.2 194.3 316.8 ;
      RECT  195.7 316.8 196.7 317.6 ;
      RECT  193.3 312.4 194.3 313.2 ;
      RECT  197.7 316.8 198.5 318.4 ;
      RECT  190.9 316.8 191.7 318.4 ;
      RECT  195.5 313.6 196.7 314.4 ;
      RECT  195.9 313.2 196.7 313.6 ;
      RECT  195.9 312.4 196.9 313.2 ;
      RECT  192.5 309.2 194.1 310.0 ;
      RECT  195.3 309.2 196.9 310.0 ;
      RECT  193.5 316.8 194.5 317.6 ;
      RECT  190.9 312.0 191.7 316.2 ;
      RECT  193.5 313.2 194.3 315.4 ;
      RECT  190.9 319.2 198.5 318.4 ;
      RECT  193.5 322.2 195.1 321.4 ;
      RECT  195.9 323.2 196.7 320.8 ;
      RECT  197.7 325.6 198.5 321.4 ;
      RECT  190.9 327.0 198.5 326.2 ;
      RECT  194.7 326.2 195.5 326.0 ;
      RECT  193.5 321.4 194.3 320.8 ;
      RECT  195.7 320.8 196.7 320.0 ;
      RECT  193.3 325.2 194.3 324.4 ;
      RECT  197.7 320.8 198.5 319.2 ;
      RECT  190.9 320.8 191.7 319.2 ;
      RECT  195.5 324.0 196.7 323.2 ;
      RECT  195.9 324.4 196.7 324.0 ;
      RECT  195.9 325.2 196.9 324.4 ;
      RECT  192.5 328.4 194.1 327.6 ;
      RECT  195.3 328.4 196.9 327.6 ;
      RECT  193.5 320.8 194.5 320.0 ;
      RECT  190.9 325.6 191.7 321.4 ;
      RECT  193.5 324.4 194.3 322.2 ;
      RECT  190.9 339.2 198.5 340.0 ;
      RECT  193.5 336.2 195.1 337.0 ;
      RECT  195.9 335.2 196.7 337.6 ;
      RECT  197.7 332.8 198.5 337.0 ;
      RECT  190.9 331.4 198.5 332.2 ;
      RECT  194.7 332.2 195.5 332.4 ;
      RECT  193.5 337.0 194.3 337.6 ;
      RECT  195.7 337.6 196.7 338.4 ;
      RECT  193.3 333.2 194.3 334.0 ;
      RECT  197.7 337.6 198.5 339.2 ;
      RECT  190.9 337.6 191.7 339.2 ;
      RECT  195.5 334.4 196.7 335.2 ;
      RECT  195.9 334.0 196.7 334.4 ;
      RECT  195.9 333.2 196.9 334.0 ;
      RECT  192.5 330.0 194.1 330.8 ;
      RECT  195.3 330.0 196.9 330.8 ;
      RECT  193.5 337.6 194.5 338.4 ;
      RECT  190.9 332.8 191.7 337.0 ;
      RECT  193.5 334.0 194.3 336.2 ;
      RECT  190.9 340.0 198.5 339.2 ;
      RECT  193.5 343.0 195.1 342.2 ;
      RECT  195.9 344.0 196.7 341.6 ;
      RECT  197.7 346.4 198.5 342.2 ;
      RECT  190.9 347.8 198.5 347.0 ;
      RECT  194.7 347.0 195.5 346.8 ;
      RECT  193.5 342.2 194.3 341.6 ;
      RECT  195.7 341.6 196.7 340.8 ;
      RECT  193.3 346.0 194.3 345.2 ;
      RECT  197.7 341.6 198.5 340.0 ;
      RECT  190.9 341.6 191.7 340.0 ;
      RECT  195.5 344.8 196.7 344.0 ;
      RECT  195.9 345.2 196.7 344.8 ;
      RECT  195.9 346.0 196.9 345.2 ;
      RECT  192.5 349.2 194.1 348.4 ;
      RECT  195.3 349.2 196.9 348.4 ;
      RECT  193.5 341.6 194.5 340.8 ;
      RECT  190.9 346.4 191.7 342.2 ;
      RECT  193.5 345.2 194.3 343.0 ;
      RECT  184.5 185.8 198.1 186.6 ;
      RECT  184.5 201.4 198.1 202.2 ;
      RECT  184.5 206.6 198.1 207.4 ;
      RECT  184.5 222.2 198.1 223.0 ;
      RECT  184.5 227.4 198.1 228.2 ;
      RECT  184.5 243.0 198.1 243.8 ;
      RECT  184.5 248.2 198.1 249.0 ;
      RECT  184.5 263.8 198.1 264.6 ;
      RECT  184.5 269.0 198.1 269.8 ;
      RECT  184.5 284.6 198.1 285.4 ;
      RECT  184.5 289.8 198.1 290.6 ;
      RECT  184.5 305.4 198.1 306.2 ;
      RECT  184.5 310.6 198.1 311.4 ;
      RECT  184.5 326.2 198.1 327.0 ;
      RECT  184.5 331.4 198.1 332.2 ;
      RECT  184.5 347.0 198.1 347.8 ;
      RECT  177.3 172.8 184.9 173.6 ;
      RECT  179.9 169.8 181.5 170.6 ;
      RECT  182.3 168.8 183.1 171.2 ;
      RECT  184.1 166.4 184.9 170.6 ;
      RECT  177.3 165.0 184.9 165.8 ;
      RECT  181.1 165.8 181.9 166.0 ;
      RECT  179.9 170.6 180.7 171.2 ;
      RECT  182.1 171.2 183.1 172.0 ;
      RECT  179.7 166.8 180.7 167.6 ;
      RECT  184.1 171.2 184.9 172.8 ;
      RECT  177.3 171.2 178.1 172.8 ;
      RECT  181.9 168.0 183.1 168.8 ;
      RECT  182.3 167.6 183.1 168.0 ;
      RECT  182.3 166.8 183.3 167.6 ;
      RECT  179.7 163.6 180.5 164.4 ;
      RECT  182.5 163.6 183.3 164.4 ;
      RECT  179.9 171.2 180.9 172.0 ;
      RECT  177.3 166.4 178.1 170.6 ;
      RECT  179.9 167.6 180.7 169.8 ;
      RECT  177.3 173.6 184.9 172.8 ;
      RECT  179.9 176.6 181.5 175.8 ;
      RECT  182.3 177.6 183.1 175.2 ;
      RECT  184.1 180.0 184.9 175.8 ;
      RECT  177.3 181.4 184.9 180.6 ;
      RECT  181.1 180.6 181.9 180.4 ;
      RECT  179.9 175.8 180.7 175.2 ;
      RECT  182.1 175.2 183.1 174.4 ;
      RECT  179.7 179.6 180.7 178.8 ;
      RECT  182.1 174.4 182.9 173.6 ;
      RECT  177.3 175.2 178.1 173.6 ;
      RECT  184.1 175.2 184.9 173.6 ;
      RECT  181.9 178.4 183.1 177.6 ;
      RECT  182.3 178.8 183.1 178.4 ;
      RECT  182.3 179.6 183.3 178.8 ;
      RECT  178.9 182.8 180.5 182.0 ;
      RECT  181.7 182.8 183.3 182.0 ;
      RECT  179.9 175.2 180.9 174.4 ;
      RECT  177.3 180.0 178.1 175.8 ;
      RECT  179.9 178.8 180.7 176.6 ;
      RECT  177.3 193.6 184.9 194.4 ;
      RECT  179.9 190.6 181.5 191.4 ;
      RECT  182.3 189.6 183.1 192.0 ;
      RECT  184.1 187.2 184.9 191.4 ;
      RECT  177.3 185.8 184.9 186.6 ;
      RECT  181.1 186.6 181.9 186.8 ;
      RECT  179.9 191.4 180.7 192.0 ;
      RECT  182.1 192.0 183.1 192.8 ;
      RECT  179.7 187.6 180.7 188.4 ;
      RECT  182.1 192.8 182.9 193.6 ;
      RECT  177.3 192.0 178.1 193.6 ;
      RECT  184.1 192.0 184.9 193.6 ;
      RECT  181.9 188.8 183.1 189.6 ;
      RECT  182.3 188.4 183.1 188.8 ;
      RECT  182.3 187.6 183.3 188.4 ;
      RECT  178.9 184.4 180.5 185.2 ;
      RECT  181.7 184.4 183.3 185.2 ;
      RECT  179.9 192.0 180.9 192.8 ;
      RECT  177.3 187.2 178.1 191.4 ;
      RECT  179.9 188.4 180.7 190.6 ;
      RECT  177.3 194.4 184.9 193.6 ;
      RECT  179.9 197.4 181.5 196.6 ;
      RECT  182.3 198.4 183.1 196.0 ;
      RECT  184.1 200.8 184.9 196.6 ;
      RECT  177.3 202.2 184.9 201.4 ;
      RECT  181.1 201.4 181.9 201.2 ;
      RECT  179.9 196.6 180.7 196.0 ;
      RECT  182.1 196.0 183.1 195.2 ;
      RECT  179.7 200.4 180.7 199.6 ;
      RECT  182.1 195.2 182.9 194.4 ;
      RECT  177.3 196.0 178.1 194.4 ;
      RECT  184.1 196.0 184.9 194.4 ;
      RECT  181.9 199.2 183.1 198.4 ;
      RECT  182.3 199.6 183.1 199.2 ;
      RECT  182.3 200.4 183.3 199.6 ;
      RECT  178.9 203.6 180.5 202.8 ;
      RECT  181.7 203.6 183.3 202.8 ;
      RECT  179.9 196.0 180.9 195.2 ;
      RECT  177.3 200.8 178.1 196.6 ;
      RECT  179.9 199.6 180.7 197.4 ;
      RECT  177.3 214.4 184.9 215.2 ;
      RECT  179.9 211.4 181.5 212.2 ;
      RECT  182.3 210.4 183.1 212.8 ;
      RECT  184.1 208.0 184.9 212.2 ;
      RECT  177.3 206.6 184.9 207.4 ;
      RECT  181.1 207.4 181.9 207.6 ;
      RECT  179.9 212.2 180.7 212.8 ;
      RECT  182.1 212.8 183.1 213.6 ;
      RECT  179.7 208.4 180.7 209.2 ;
      RECT  182.1 213.6 182.9 214.4 ;
      RECT  177.3 212.8 178.1 214.4 ;
      RECT  184.1 212.8 184.9 214.4 ;
      RECT  181.9 209.6 183.1 210.4 ;
      RECT  182.3 209.2 183.1 209.6 ;
      RECT  182.3 208.4 183.3 209.2 ;
      RECT  178.9 205.2 180.5 206.0 ;
      RECT  181.7 205.2 183.3 206.0 ;
      RECT  179.9 212.8 180.9 213.6 ;
      RECT  177.3 208.0 178.1 212.2 ;
      RECT  179.9 209.2 180.7 211.4 ;
      RECT  177.3 215.2 184.9 214.4 ;
      RECT  179.9 218.2 181.5 217.4 ;
      RECT  182.3 219.2 183.1 216.8 ;
      RECT  184.1 221.6 184.9 217.4 ;
      RECT  177.3 223.0 184.9 222.2 ;
      RECT  181.1 222.2 181.9 222.0 ;
      RECT  179.9 217.4 180.7 216.8 ;
      RECT  182.1 216.8 183.1 216.0 ;
      RECT  179.7 221.2 180.7 220.4 ;
      RECT  182.1 216.0 182.9 215.2 ;
      RECT  177.3 216.8 178.1 215.2 ;
      RECT  184.1 216.8 184.9 215.2 ;
      RECT  181.9 220.0 183.1 219.2 ;
      RECT  182.3 220.4 183.1 220.0 ;
      RECT  182.3 221.2 183.3 220.4 ;
      RECT  178.9 224.4 180.5 223.6 ;
      RECT  181.7 224.4 183.3 223.6 ;
      RECT  179.9 216.8 180.9 216.0 ;
      RECT  177.3 221.6 178.1 217.4 ;
      RECT  179.9 220.4 180.7 218.2 ;
      RECT  177.3 235.2 184.9 236.0 ;
      RECT  179.9 232.2 181.5 233.0 ;
      RECT  182.3 231.2 183.1 233.6 ;
      RECT  184.1 228.8 184.9 233.0 ;
      RECT  177.3 227.4 184.9 228.2 ;
      RECT  181.1 228.2 181.9 228.4 ;
      RECT  179.9 233.0 180.7 233.6 ;
      RECT  182.1 233.6 183.1 234.4 ;
      RECT  179.7 229.2 180.7 230.0 ;
      RECT  182.1 234.4 182.9 235.2 ;
      RECT  177.3 233.6 178.1 235.2 ;
      RECT  184.1 233.6 184.9 235.2 ;
      RECT  181.9 230.4 183.1 231.2 ;
      RECT  182.3 230.0 183.1 230.4 ;
      RECT  182.3 229.2 183.3 230.0 ;
      RECT  178.9 226.0 180.5 226.8 ;
      RECT  181.7 226.0 183.3 226.8 ;
      RECT  179.9 233.6 180.9 234.4 ;
      RECT  177.3 228.8 178.1 233.0 ;
      RECT  179.9 230.0 180.7 232.2 ;
      RECT  177.3 236.0 184.9 235.2 ;
      RECT  179.9 239.0 181.5 238.2 ;
      RECT  182.3 240.0 183.1 237.6 ;
      RECT  184.1 242.4 184.9 238.2 ;
      RECT  177.3 243.8 184.9 243.0 ;
      RECT  181.1 243.0 181.9 242.8 ;
      RECT  179.9 238.2 180.7 237.6 ;
      RECT  182.1 237.6 183.1 236.8 ;
      RECT  179.7 242.0 180.7 241.2 ;
      RECT  182.1 236.8 182.9 236.0 ;
      RECT  177.3 237.6 178.1 236.0 ;
      RECT  184.1 237.6 184.9 236.0 ;
      RECT  181.9 240.8 183.1 240.0 ;
      RECT  182.3 241.2 183.1 240.8 ;
      RECT  182.3 242.0 183.3 241.2 ;
      RECT  178.9 245.2 180.5 244.4 ;
      RECT  181.7 245.2 183.3 244.4 ;
      RECT  179.9 237.6 180.9 236.8 ;
      RECT  177.3 242.4 178.1 238.2 ;
      RECT  179.9 241.2 180.7 239.0 ;
      RECT  177.3 256.0 184.9 256.8 ;
      RECT  179.9 253.0 181.5 253.8 ;
      RECT  182.3 252.0 183.1 254.4 ;
      RECT  184.1 249.6 184.9 253.8 ;
      RECT  177.3 248.2 184.9 249.0 ;
      RECT  181.1 249.0 181.9 249.2 ;
      RECT  179.9 253.8 180.7 254.4 ;
      RECT  182.1 254.4 183.1 255.2 ;
      RECT  179.7 250.0 180.7 250.8 ;
      RECT  182.1 255.2 182.9 256.0 ;
      RECT  177.3 254.4 178.1 256.0 ;
      RECT  184.1 254.4 184.9 256.0 ;
      RECT  181.9 251.2 183.1 252.0 ;
      RECT  182.3 250.8 183.1 251.2 ;
      RECT  182.3 250.0 183.3 250.8 ;
      RECT  178.9 246.8 180.5 247.6 ;
      RECT  181.7 246.8 183.3 247.6 ;
      RECT  179.9 254.4 180.9 255.2 ;
      RECT  177.3 249.6 178.1 253.8 ;
      RECT  179.9 250.8 180.7 253.0 ;
      RECT  177.3 256.8 184.9 256.0 ;
      RECT  179.9 259.8 181.5 259.0 ;
      RECT  182.3 260.8 183.1 258.4 ;
      RECT  184.1 263.2 184.9 259.0 ;
      RECT  177.3 264.6 184.9 263.8 ;
      RECT  181.1 263.8 181.9 263.6 ;
      RECT  179.9 259.0 180.7 258.4 ;
      RECT  182.1 258.4 183.1 257.6 ;
      RECT  179.7 262.8 180.7 262.0 ;
      RECT  182.1 257.6 182.9 256.8 ;
      RECT  177.3 258.4 178.1 256.8 ;
      RECT  184.1 258.4 184.9 256.8 ;
      RECT  181.9 261.6 183.1 260.8 ;
      RECT  182.3 262.0 183.1 261.6 ;
      RECT  182.3 262.8 183.3 262.0 ;
      RECT  178.9 266.0 180.5 265.2 ;
      RECT  181.7 266.0 183.3 265.2 ;
      RECT  179.9 258.4 180.9 257.6 ;
      RECT  177.3 263.2 178.1 259.0 ;
      RECT  179.9 262.0 180.7 259.8 ;
      RECT  177.3 276.8 184.9 277.6 ;
      RECT  179.9 273.8 181.5 274.6 ;
      RECT  182.3 272.8 183.1 275.2 ;
      RECT  184.1 270.4 184.9 274.6 ;
      RECT  177.3 269.0 184.9 269.8 ;
      RECT  181.1 269.8 181.9 270.0 ;
      RECT  179.9 274.6 180.7 275.2 ;
      RECT  182.1 275.2 183.1 276.0 ;
      RECT  179.7 270.8 180.7 271.6 ;
      RECT  182.1 276.0 182.9 276.8 ;
      RECT  177.3 275.2 178.1 276.8 ;
      RECT  184.1 275.2 184.9 276.8 ;
      RECT  181.9 272.0 183.1 272.8 ;
      RECT  182.3 271.6 183.1 272.0 ;
      RECT  182.3 270.8 183.3 271.6 ;
      RECT  178.9 267.6 180.5 268.4 ;
      RECT  181.7 267.6 183.3 268.4 ;
      RECT  179.9 275.2 180.9 276.0 ;
      RECT  177.3 270.4 178.1 274.6 ;
      RECT  179.9 271.6 180.7 273.8 ;
      RECT  177.3 277.6 184.9 276.8 ;
      RECT  179.9 280.6 181.5 279.8 ;
      RECT  182.3 281.6 183.1 279.2 ;
      RECT  184.1 284.0 184.9 279.8 ;
      RECT  177.3 285.4 184.9 284.6 ;
      RECT  181.1 284.6 181.9 284.4 ;
      RECT  179.9 279.8 180.7 279.2 ;
      RECT  182.1 279.2 183.1 278.4 ;
      RECT  179.7 283.6 180.7 282.8 ;
      RECT  182.1 278.4 182.9 277.6 ;
      RECT  177.3 279.2 178.1 277.6 ;
      RECT  184.1 279.2 184.9 277.6 ;
      RECT  181.9 282.4 183.1 281.6 ;
      RECT  182.3 282.8 183.1 282.4 ;
      RECT  182.3 283.6 183.3 282.8 ;
      RECT  178.9 286.8 180.5 286.0 ;
      RECT  181.7 286.8 183.3 286.0 ;
      RECT  179.9 279.2 180.9 278.4 ;
      RECT  177.3 284.0 178.1 279.8 ;
      RECT  179.9 282.8 180.7 280.6 ;
      RECT  177.3 297.6 184.9 298.4 ;
      RECT  179.9 294.6 181.5 295.4 ;
      RECT  182.3 293.6 183.1 296.0 ;
      RECT  184.1 291.2 184.9 295.4 ;
      RECT  177.3 289.8 184.9 290.6 ;
      RECT  181.1 290.6 181.9 290.8 ;
      RECT  179.9 295.4 180.7 296.0 ;
      RECT  182.1 296.0 183.1 296.8 ;
      RECT  179.7 291.6 180.7 292.4 ;
      RECT  182.1 296.8 182.9 297.6 ;
      RECT  177.3 296.0 178.1 297.6 ;
      RECT  184.1 296.0 184.9 297.6 ;
      RECT  181.9 292.8 183.1 293.6 ;
      RECT  182.3 292.4 183.1 292.8 ;
      RECT  182.3 291.6 183.3 292.4 ;
      RECT  178.9 288.4 180.5 289.2 ;
      RECT  181.7 288.4 183.3 289.2 ;
      RECT  179.9 296.0 180.9 296.8 ;
      RECT  177.3 291.2 178.1 295.4 ;
      RECT  179.9 292.4 180.7 294.6 ;
      RECT  177.3 298.4 184.9 297.6 ;
      RECT  179.9 301.4 181.5 300.6 ;
      RECT  182.3 302.4 183.1 300.0 ;
      RECT  184.1 304.8 184.9 300.6 ;
      RECT  177.3 306.2 184.9 305.4 ;
      RECT  181.1 305.4 181.9 305.2 ;
      RECT  179.9 300.6 180.7 300.0 ;
      RECT  182.1 300.0 183.1 299.2 ;
      RECT  179.7 304.4 180.7 303.6 ;
      RECT  182.1 299.2 182.9 298.4 ;
      RECT  177.3 300.0 178.1 298.4 ;
      RECT  184.1 300.0 184.9 298.4 ;
      RECT  181.9 303.2 183.1 302.4 ;
      RECT  182.3 303.6 183.1 303.2 ;
      RECT  182.3 304.4 183.3 303.6 ;
      RECT  178.9 307.6 180.5 306.8 ;
      RECT  181.7 307.6 183.3 306.8 ;
      RECT  179.9 300.0 180.9 299.2 ;
      RECT  177.3 304.8 178.1 300.6 ;
      RECT  179.9 303.6 180.7 301.4 ;
      RECT  177.3 318.4 184.9 319.2 ;
      RECT  179.9 315.4 181.5 316.2 ;
      RECT  182.3 314.4 183.1 316.8 ;
      RECT  184.1 312.0 184.9 316.2 ;
      RECT  177.3 310.6 184.9 311.4 ;
      RECT  181.1 311.4 181.9 311.6 ;
      RECT  179.9 316.2 180.7 316.8 ;
      RECT  182.1 316.8 183.1 317.6 ;
      RECT  179.7 312.4 180.7 313.2 ;
      RECT  182.1 317.6 182.9 318.4 ;
      RECT  177.3 316.8 178.1 318.4 ;
      RECT  184.1 316.8 184.9 318.4 ;
      RECT  181.9 313.6 183.1 314.4 ;
      RECT  182.3 313.2 183.1 313.6 ;
      RECT  182.3 312.4 183.3 313.2 ;
      RECT  178.9 309.2 180.5 310.0 ;
      RECT  181.7 309.2 183.3 310.0 ;
      RECT  179.9 316.8 180.9 317.6 ;
      RECT  177.3 312.0 178.1 316.2 ;
      RECT  179.9 313.2 180.7 315.4 ;
      RECT  177.3 319.2 184.9 318.4 ;
      RECT  179.9 322.2 181.5 321.4 ;
      RECT  182.3 323.2 183.1 320.8 ;
      RECT  184.1 325.6 184.9 321.4 ;
      RECT  177.3 327.0 184.9 326.2 ;
      RECT  181.1 326.2 181.9 326.0 ;
      RECT  179.9 321.4 180.7 320.8 ;
      RECT  182.1 320.8 183.1 320.0 ;
      RECT  179.7 325.2 180.7 324.4 ;
      RECT  182.1 320.0 182.9 319.2 ;
      RECT  177.3 320.8 178.1 319.2 ;
      RECT  184.1 320.8 184.9 319.2 ;
      RECT  181.9 324.0 183.1 323.2 ;
      RECT  182.3 324.4 183.1 324.0 ;
      RECT  182.3 325.2 183.3 324.4 ;
      RECT  178.9 328.4 180.5 327.6 ;
      RECT  181.7 328.4 183.3 327.6 ;
      RECT  179.9 320.8 180.9 320.0 ;
      RECT  177.3 325.6 178.1 321.4 ;
      RECT  179.9 324.4 180.7 322.2 ;
      RECT  177.3 339.2 184.9 340.0 ;
      RECT  179.9 336.2 181.5 337.0 ;
      RECT  182.3 335.2 183.1 337.6 ;
      RECT  184.1 332.8 184.9 337.0 ;
      RECT  177.3 331.4 184.9 332.2 ;
      RECT  181.1 332.2 181.9 332.4 ;
      RECT  179.9 337.0 180.7 337.6 ;
      RECT  182.1 337.6 183.1 338.4 ;
      RECT  179.7 333.2 180.7 334.0 ;
      RECT  182.1 338.4 182.9 339.2 ;
      RECT  177.3 337.6 178.1 339.2 ;
      RECT  184.1 337.6 184.9 339.2 ;
      RECT  181.9 334.4 183.1 335.2 ;
      RECT  182.3 334.0 183.1 334.4 ;
      RECT  182.3 333.2 183.3 334.0 ;
      RECT  178.9 330.0 180.5 330.8 ;
      RECT  181.7 330.0 183.3 330.8 ;
      RECT  179.9 337.6 180.9 338.4 ;
      RECT  177.3 332.8 178.1 337.0 ;
      RECT  179.9 334.0 180.7 336.2 ;
      RECT  177.3 340.0 184.9 339.2 ;
      RECT  179.9 343.0 181.5 342.2 ;
      RECT  182.3 344.0 183.1 341.6 ;
      RECT  184.1 346.4 184.9 342.2 ;
      RECT  177.3 347.8 184.9 347.0 ;
      RECT  181.1 347.0 181.9 346.8 ;
      RECT  179.9 342.2 180.7 341.6 ;
      RECT  182.1 341.6 183.1 340.8 ;
      RECT  179.7 346.0 180.7 345.2 ;
      RECT  182.1 340.8 182.9 340.0 ;
      RECT  177.3 341.6 178.1 340.0 ;
      RECT  184.1 341.6 184.9 340.0 ;
      RECT  181.9 344.8 183.1 344.0 ;
      RECT  182.3 345.2 183.1 344.8 ;
      RECT  182.3 346.0 183.3 345.2 ;
      RECT  178.9 349.2 180.5 348.4 ;
      RECT  181.7 349.2 183.3 348.4 ;
      RECT  179.9 341.6 180.9 340.8 ;
      RECT  177.3 346.4 178.1 342.2 ;
      RECT  179.9 345.2 180.7 343.0 ;
      RECT  177.3 360.0 184.9 360.8 ;
      RECT  179.9 357.0 181.5 357.8 ;
      RECT  182.3 356.0 183.1 358.4 ;
      RECT  184.1 353.6 184.9 357.8 ;
      RECT  177.3 352.2 184.9 353.0 ;
      RECT  181.1 353.0 181.9 353.2 ;
      RECT  179.9 357.8 180.7 358.4 ;
      RECT  182.1 358.4 183.1 359.2 ;
      RECT  179.7 354.0 180.7 354.8 ;
      RECT  184.1 358.4 184.9 360.0 ;
      RECT  177.3 358.4 178.1 360.0 ;
      RECT  181.9 355.2 183.1 356.0 ;
      RECT  182.3 354.8 183.1 355.2 ;
      RECT  182.3 354.0 183.3 354.8 ;
      RECT  179.7 350.8 180.5 351.6 ;
      RECT  182.5 350.8 183.3 351.6 ;
      RECT  179.9 358.4 180.9 359.2 ;
      RECT  177.3 353.6 178.1 357.8 ;
      RECT  179.9 354.8 180.7 357.0 ;
      RECT  177.7 165.0 184.5 165.8 ;
      RECT  177.7 180.6 184.5 181.4 ;
      RECT  177.7 185.8 184.5 186.6 ;
      RECT  177.7 201.4 184.5 202.2 ;
      RECT  177.7 206.6 184.5 207.4 ;
      RECT  177.7 222.2 184.5 223.0 ;
      RECT  177.7 227.4 184.5 228.2 ;
      RECT  177.7 243.0 184.5 243.8 ;
      RECT  177.7 248.2 184.5 249.0 ;
      RECT  177.7 263.8 184.5 264.6 ;
      RECT  177.7 269.0 184.5 269.8 ;
      RECT  177.7 284.6 184.5 285.4 ;
      RECT  177.7 289.8 184.5 290.6 ;
      RECT  177.7 305.4 184.5 306.2 ;
      RECT  177.7 310.6 184.5 311.4 ;
      RECT  177.7 326.2 184.5 327.0 ;
      RECT  177.7 331.4 184.5 332.2 ;
      RECT  177.7 347.0 184.5 347.8 ;
      RECT  177.7 352.2 184.5 353.0 ;
      RECT  184.1 173.6 191.7 172.8 ;
      RECT  186.7 176.6 188.3 175.8 ;
      RECT  189.1 177.6 189.9 175.2 ;
      RECT  190.9 180.0 191.7 175.8 ;
      RECT  184.1 181.4 191.7 180.6 ;
      RECT  187.9 180.6 188.7 180.4 ;
      RECT  186.7 175.8 187.5 175.2 ;
      RECT  188.9 175.2 189.9 174.4 ;
      RECT  186.5 179.6 187.5 178.8 ;
      RECT  190.9 175.2 191.7 173.6 ;
      RECT  184.1 175.2 184.9 173.6 ;
      RECT  188.7 178.4 189.9 177.6 ;
      RECT  189.1 178.8 189.9 178.4 ;
      RECT  189.1 179.6 190.1 178.8 ;
      RECT  186.5 182.8 187.3 182.0 ;
      RECT  189.3 182.8 190.1 182.0 ;
      RECT  186.7 175.2 187.7 174.4 ;
      RECT  184.1 180.0 184.9 175.8 ;
      RECT  186.7 178.8 187.5 176.6 ;
      RECT  190.9 173.6 198.5 172.8 ;
      RECT  193.5 176.6 195.1 175.8 ;
      RECT  195.9 177.6 196.7 175.2 ;
      RECT  197.7 180.0 198.5 175.8 ;
      RECT  190.9 181.4 198.5 180.6 ;
      RECT  194.7 180.6 195.5 180.4 ;
      RECT  193.5 175.8 194.3 175.2 ;
      RECT  195.7 175.2 196.7 174.4 ;
      RECT  193.3 179.6 194.3 178.8 ;
      RECT  197.7 175.2 198.5 173.6 ;
      RECT  190.9 175.2 191.7 173.6 ;
      RECT  195.5 178.4 196.7 177.6 ;
      RECT  195.9 178.8 196.7 178.4 ;
      RECT  195.9 179.6 196.9 178.8 ;
      RECT  193.3 182.8 194.1 182.0 ;
      RECT  196.1 182.8 196.9 182.0 ;
      RECT  193.5 175.2 194.5 174.4 ;
      RECT  190.9 180.0 191.7 175.8 ;
      RECT  193.5 178.8 194.3 176.6 ;
      RECT  184.5 181.4 198.1 180.6 ;
      RECT  184.1 172.8 191.7 173.6 ;
      RECT  186.7 169.8 188.3 170.6 ;
      RECT  189.1 168.8 189.9 171.2 ;
      RECT  190.9 166.4 191.7 170.6 ;
      RECT  184.1 165.0 191.7 165.8 ;
      RECT  187.9 165.8 188.7 166.0 ;
      RECT  186.7 170.6 187.5 171.2 ;
      RECT  188.9 171.2 189.9 172.0 ;
      RECT  186.5 166.8 187.5 167.6 ;
      RECT  190.9 171.2 191.7 172.8 ;
      RECT  184.1 171.2 184.9 172.8 ;
      RECT  188.7 168.0 189.9 168.8 ;
      RECT  189.1 167.6 189.9 168.0 ;
      RECT  189.1 166.8 190.1 167.6 ;
      RECT  186.5 163.6 187.3 164.4 ;
      RECT  189.3 163.6 190.1 164.4 ;
      RECT  186.7 171.2 187.7 172.0 ;
      RECT  184.1 166.4 184.9 170.6 ;
      RECT  186.7 167.6 187.5 169.8 ;
      RECT  190.9 172.8 198.5 173.6 ;
      RECT  193.5 169.8 195.1 170.6 ;
      RECT  195.9 168.8 196.7 171.2 ;
      RECT  197.7 166.4 198.5 170.6 ;
      RECT  190.9 165.0 198.5 165.8 ;
      RECT  194.7 165.8 195.5 166.0 ;
      RECT  193.5 170.6 194.3 171.2 ;
      RECT  195.7 171.2 196.7 172.0 ;
      RECT  193.3 166.8 194.3 167.6 ;
      RECT  197.7 171.2 198.5 172.8 ;
      RECT  190.9 171.2 191.7 172.8 ;
      RECT  195.5 168.0 196.7 168.8 ;
      RECT  195.9 167.6 196.7 168.0 ;
      RECT  195.9 166.8 196.9 167.6 ;
      RECT  193.3 163.6 194.1 164.4 ;
      RECT  196.1 163.6 196.9 164.4 ;
      RECT  193.5 171.2 194.5 172.0 ;
      RECT  190.9 166.4 191.7 170.6 ;
      RECT  193.5 167.6 194.3 169.8 ;
      RECT  184.5 165.0 198.1 165.8 ;
      RECT  184.1 360.0 191.7 360.8 ;
      RECT  186.7 357.0 188.3 357.8 ;
      RECT  189.1 356.0 189.9 358.4 ;
      RECT  190.9 353.6 191.7 357.8 ;
      RECT  184.1 352.2 191.7 353.0 ;
      RECT  187.9 353.0 188.7 353.2 ;
      RECT  186.7 357.8 187.5 358.4 ;
      RECT  188.9 358.4 189.9 359.2 ;
      RECT  186.5 354.0 187.5 354.8 ;
      RECT  190.9 358.4 191.7 360.0 ;
      RECT  184.1 358.4 184.9 360.0 ;
      RECT  188.7 355.2 189.9 356.0 ;
      RECT  189.1 354.8 189.9 355.2 ;
      RECT  189.1 354.0 190.1 354.8 ;
      RECT  186.5 350.8 187.3 351.6 ;
      RECT  189.3 350.8 190.1 351.6 ;
      RECT  186.7 358.4 187.7 359.2 ;
      RECT  184.1 353.6 184.9 357.8 ;
      RECT  186.7 354.8 187.5 357.0 ;
      RECT  190.9 360.0 198.5 360.8 ;
      RECT  193.5 357.0 195.1 357.8 ;
      RECT  195.9 356.0 196.7 358.4 ;
      RECT  197.7 353.6 198.5 357.8 ;
      RECT  190.9 352.2 198.5 353.0 ;
      RECT  194.7 353.0 195.5 353.2 ;
      RECT  193.5 357.8 194.3 358.4 ;
      RECT  195.7 358.4 196.7 359.2 ;
      RECT  193.3 354.0 194.3 354.8 ;
      RECT  197.7 358.4 198.5 360.0 ;
      RECT  190.9 358.4 191.7 360.0 ;
      RECT  195.5 355.2 196.7 356.0 ;
      RECT  195.9 354.8 196.7 355.2 ;
      RECT  195.9 354.0 196.9 354.8 ;
      RECT  193.3 350.8 194.1 351.6 ;
      RECT  196.1 350.8 196.9 351.6 ;
      RECT  193.5 358.4 194.5 359.2 ;
      RECT  190.9 353.6 191.7 357.8 ;
      RECT  193.5 354.8 194.3 357.0 ;
      RECT  184.5 352.2 198.1 353.0 ;
      RECT  170.5 172.8 178.1 173.6 ;
      RECT  173.1 169.8 174.7 170.6 ;
      RECT  175.5 168.8 176.3 171.2 ;
      RECT  177.3 166.4 178.1 170.6 ;
      RECT  170.5 165.0 178.1 165.8 ;
      RECT  174.3 165.8 175.1 166.0 ;
      RECT  173.1 170.6 173.9 171.2 ;
      RECT  175.3 171.2 176.3 172.0 ;
      RECT  172.9 166.8 173.9 167.6 ;
      RECT  177.3 171.2 178.1 172.8 ;
      RECT  170.5 171.2 171.3 172.8 ;
      RECT  175.1 168.0 176.3 168.8 ;
      RECT  175.5 167.6 176.3 168.0 ;
      RECT  175.5 166.8 176.5 167.6 ;
      RECT  172.9 163.6 173.7 164.4 ;
      RECT  175.7 163.6 176.5 164.4 ;
      RECT  173.1 171.2 174.1 172.0 ;
      RECT  170.5 166.4 171.3 170.6 ;
      RECT  173.1 167.6 173.9 169.8 ;
      RECT  170.5 173.6 178.1 172.8 ;
      RECT  173.1 176.6 174.7 175.8 ;
      RECT  175.5 177.6 176.3 175.2 ;
      RECT  177.3 180.0 178.1 175.8 ;
      RECT  170.5 181.4 178.1 180.6 ;
      RECT  174.3 180.6 175.1 180.4 ;
      RECT  173.1 175.8 173.9 175.2 ;
      RECT  175.3 175.2 176.3 174.4 ;
      RECT  172.9 179.6 173.9 178.8 ;
      RECT  177.3 175.2 178.1 173.6 ;
      RECT  170.5 175.2 171.3 173.6 ;
      RECT  175.1 178.4 176.3 177.6 ;
      RECT  175.5 178.8 176.3 178.4 ;
      RECT  175.5 179.6 176.5 178.8 ;
      RECT  172.9 182.8 173.7 182.0 ;
      RECT  175.7 182.8 176.5 182.0 ;
      RECT  173.1 175.2 174.1 174.4 ;
      RECT  170.5 180.0 171.3 175.8 ;
      RECT  173.1 178.8 173.9 176.6 ;
      RECT  170.5 193.6 178.1 194.4 ;
      RECT  173.1 190.6 174.7 191.4 ;
      RECT  175.5 189.6 176.3 192.0 ;
      RECT  177.3 187.2 178.1 191.4 ;
      RECT  170.5 185.8 178.1 186.6 ;
      RECT  174.3 186.6 175.1 186.8 ;
      RECT  173.1 191.4 173.9 192.0 ;
      RECT  175.3 192.0 176.3 192.8 ;
      RECT  172.9 187.6 173.9 188.4 ;
      RECT  177.3 192.0 178.1 193.6 ;
      RECT  170.5 192.0 171.3 193.6 ;
      RECT  175.1 188.8 176.3 189.6 ;
      RECT  175.5 188.4 176.3 188.8 ;
      RECT  175.5 187.6 176.5 188.4 ;
      RECT  172.9 184.4 173.7 185.2 ;
      RECT  175.7 184.4 176.5 185.2 ;
      RECT  173.1 192.0 174.1 192.8 ;
      RECT  170.5 187.2 171.3 191.4 ;
      RECT  173.1 188.4 173.9 190.6 ;
      RECT  170.5 194.4 178.1 193.6 ;
      RECT  173.1 197.4 174.7 196.6 ;
      RECT  175.5 198.4 176.3 196.0 ;
      RECT  177.3 200.8 178.1 196.6 ;
      RECT  170.5 202.2 178.1 201.4 ;
      RECT  174.3 201.4 175.1 201.2 ;
      RECT  173.1 196.6 173.9 196.0 ;
      RECT  175.3 196.0 176.3 195.2 ;
      RECT  172.9 200.4 173.9 199.6 ;
      RECT  177.3 196.0 178.1 194.4 ;
      RECT  170.5 196.0 171.3 194.4 ;
      RECT  175.1 199.2 176.3 198.4 ;
      RECT  175.5 199.6 176.3 199.2 ;
      RECT  175.5 200.4 176.5 199.6 ;
      RECT  172.9 203.6 173.7 202.8 ;
      RECT  175.7 203.6 176.5 202.8 ;
      RECT  173.1 196.0 174.1 195.2 ;
      RECT  170.5 200.8 171.3 196.6 ;
      RECT  173.1 199.6 173.9 197.4 ;
      RECT  170.5 214.4 178.1 215.2 ;
      RECT  173.1 211.4 174.7 212.2 ;
      RECT  175.5 210.4 176.3 212.8 ;
      RECT  177.3 208.0 178.1 212.2 ;
      RECT  170.5 206.6 178.1 207.4 ;
      RECT  174.3 207.4 175.1 207.6 ;
      RECT  173.1 212.2 173.9 212.8 ;
      RECT  175.3 212.8 176.3 213.6 ;
      RECT  172.9 208.4 173.9 209.2 ;
      RECT  177.3 212.8 178.1 214.4 ;
      RECT  170.5 212.8 171.3 214.4 ;
      RECT  175.1 209.6 176.3 210.4 ;
      RECT  175.5 209.2 176.3 209.6 ;
      RECT  175.5 208.4 176.5 209.2 ;
      RECT  172.9 205.2 173.7 206.0 ;
      RECT  175.7 205.2 176.5 206.0 ;
      RECT  173.1 212.8 174.1 213.6 ;
      RECT  170.5 208.0 171.3 212.2 ;
      RECT  173.1 209.2 173.9 211.4 ;
      RECT  170.5 215.2 178.1 214.4 ;
      RECT  173.1 218.2 174.7 217.4 ;
      RECT  175.5 219.2 176.3 216.8 ;
      RECT  177.3 221.6 178.1 217.4 ;
      RECT  170.5 223.0 178.1 222.2 ;
      RECT  174.3 222.2 175.1 222.0 ;
      RECT  173.1 217.4 173.9 216.8 ;
      RECT  175.3 216.8 176.3 216.0 ;
      RECT  172.9 221.2 173.9 220.4 ;
      RECT  177.3 216.8 178.1 215.2 ;
      RECT  170.5 216.8 171.3 215.2 ;
      RECT  175.1 220.0 176.3 219.2 ;
      RECT  175.5 220.4 176.3 220.0 ;
      RECT  175.5 221.2 176.5 220.4 ;
      RECT  172.9 224.4 173.7 223.6 ;
      RECT  175.7 224.4 176.5 223.6 ;
      RECT  173.1 216.8 174.1 216.0 ;
      RECT  170.5 221.6 171.3 217.4 ;
      RECT  173.1 220.4 173.9 218.2 ;
      RECT  170.5 235.2 178.1 236.0 ;
      RECT  173.1 232.2 174.7 233.0 ;
      RECT  175.5 231.2 176.3 233.6 ;
      RECT  177.3 228.8 178.1 233.0 ;
      RECT  170.5 227.4 178.1 228.2 ;
      RECT  174.3 228.2 175.1 228.4 ;
      RECT  173.1 233.0 173.9 233.6 ;
      RECT  175.3 233.6 176.3 234.4 ;
      RECT  172.9 229.2 173.9 230.0 ;
      RECT  177.3 233.6 178.1 235.2 ;
      RECT  170.5 233.6 171.3 235.2 ;
      RECT  175.1 230.4 176.3 231.2 ;
      RECT  175.5 230.0 176.3 230.4 ;
      RECT  175.5 229.2 176.5 230.0 ;
      RECT  172.9 226.0 173.7 226.8 ;
      RECT  175.7 226.0 176.5 226.8 ;
      RECT  173.1 233.6 174.1 234.4 ;
      RECT  170.5 228.8 171.3 233.0 ;
      RECT  173.1 230.0 173.9 232.2 ;
      RECT  170.5 236.0 178.1 235.2 ;
      RECT  173.1 239.0 174.7 238.2 ;
      RECT  175.5 240.0 176.3 237.6 ;
      RECT  177.3 242.4 178.1 238.2 ;
      RECT  170.5 243.8 178.1 243.0 ;
      RECT  174.3 243.0 175.1 242.8 ;
      RECT  173.1 238.2 173.9 237.6 ;
      RECT  175.3 237.6 176.3 236.8 ;
      RECT  172.9 242.0 173.9 241.2 ;
      RECT  177.3 237.6 178.1 236.0 ;
      RECT  170.5 237.6 171.3 236.0 ;
      RECT  175.1 240.8 176.3 240.0 ;
      RECT  175.5 241.2 176.3 240.8 ;
      RECT  175.5 242.0 176.5 241.2 ;
      RECT  172.9 245.2 173.7 244.4 ;
      RECT  175.7 245.2 176.5 244.4 ;
      RECT  173.1 237.6 174.1 236.8 ;
      RECT  170.5 242.4 171.3 238.2 ;
      RECT  173.1 241.2 173.9 239.0 ;
      RECT  170.5 256.0 178.1 256.8 ;
      RECT  173.1 253.0 174.7 253.8 ;
      RECT  175.5 252.0 176.3 254.4 ;
      RECT  177.3 249.6 178.1 253.8 ;
      RECT  170.5 248.2 178.1 249.0 ;
      RECT  174.3 249.0 175.1 249.2 ;
      RECT  173.1 253.8 173.9 254.4 ;
      RECT  175.3 254.4 176.3 255.2 ;
      RECT  172.9 250.0 173.9 250.8 ;
      RECT  177.3 254.4 178.1 256.0 ;
      RECT  170.5 254.4 171.3 256.0 ;
      RECT  175.1 251.2 176.3 252.0 ;
      RECT  175.5 250.8 176.3 251.2 ;
      RECT  175.5 250.0 176.5 250.8 ;
      RECT  172.9 246.8 173.7 247.6 ;
      RECT  175.7 246.8 176.5 247.6 ;
      RECT  173.1 254.4 174.1 255.2 ;
      RECT  170.5 249.6 171.3 253.8 ;
      RECT  173.1 250.8 173.9 253.0 ;
      RECT  170.5 256.8 178.1 256.0 ;
      RECT  173.1 259.8 174.7 259.0 ;
      RECT  175.5 260.8 176.3 258.4 ;
      RECT  177.3 263.2 178.1 259.0 ;
      RECT  170.5 264.6 178.1 263.8 ;
      RECT  174.3 263.8 175.1 263.6 ;
      RECT  173.1 259.0 173.9 258.4 ;
      RECT  175.3 258.4 176.3 257.6 ;
      RECT  172.9 262.8 173.9 262.0 ;
      RECT  177.3 258.4 178.1 256.8 ;
      RECT  170.5 258.4 171.3 256.8 ;
      RECT  175.1 261.6 176.3 260.8 ;
      RECT  175.5 262.0 176.3 261.6 ;
      RECT  175.5 262.8 176.5 262.0 ;
      RECT  172.9 266.0 173.7 265.2 ;
      RECT  175.7 266.0 176.5 265.2 ;
      RECT  173.1 258.4 174.1 257.6 ;
      RECT  170.5 263.2 171.3 259.0 ;
      RECT  173.1 262.0 173.9 259.8 ;
      RECT  170.5 276.8 178.1 277.6 ;
      RECT  173.1 273.8 174.7 274.6 ;
      RECT  175.5 272.8 176.3 275.2 ;
      RECT  177.3 270.4 178.1 274.6 ;
      RECT  170.5 269.0 178.1 269.8 ;
      RECT  174.3 269.8 175.1 270.0 ;
      RECT  173.1 274.6 173.9 275.2 ;
      RECT  175.3 275.2 176.3 276.0 ;
      RECT  172.9 270.8 173.9 271.6 ;
      RECT  177.3 275.2 178.1 276.8 ;
      RECT  170.5 275.2 171.3 276.8 ;
      RECT  175.1 272.0 176.3 272.8 ;
      RECT  175.5 271.6 176.3 272.0 ;
      RECT  175.5 270.8 176.5 271.6 ;
      RECT  172.9 267.6 173.7 268.4 ;
      RECT  175.7 267.6 176.5 268.4 ;
      RECT  173.1 275.2 174.1 276.0 ;
      RECT  170.5 270.4 171.3 274.6 ;
      RECT  173.1 271.6 173.9 273.8 ;
      RECT  170.5 277.6 178.1 276.8 ;
      RECT  173.1 280.6 174.7 279.8 ;
      RECT  175.5 281.6 176.3 279.2 ;
      RECT  177.3 284.0 178.1 279.8 ;
      RECT  170.5 285.4 178.1 284.6 ;
      RECT  174.3 284.6 175.1 284.4 ;
      RECT  173.1 279.8 173.9 279.2 ;
      RECT  175.3 279.2 176.3 278.4 ;
      RECT  172.9 283.6 173.9 282.8 ;
      RECT  177.3 279.2 178.1 277.6 ;
      RECT  170.5 279.2 171.3 277.6 ;
      RECT  175.1 282.4 176.3 281.6 ;
      RECT  175.5 282.8 176.3 282.4 ;
      RECT  175.5 283.6 176.5 282.8 ;
      RECT  172.9 286.8 173.7 286.0 ;
      RECT  175.7 286.8 176.5 286.0 ;
      RECT  173.1 279.2 174.1 278.4 ;
      RECT  170.5 284.0 171.3 279.8 ;
      RECT  173.1 282.8 173.9 280.6 ;
      RECT  170.5 297.6 178.1 298.4 ;
      RECT  173.1 294.6 174.7 295.4 ;
      RECT  175.5 293.6 176.3 296.0 ;
      RECT  177.3 291.2 178.1 295.4 ;
      RECT  170.5 289.8 178.1 290.6 ;
      RECT  174.3 290.6 175.1 290.8 ;
      RECT  173.1 295.4 173.9 296.0 ;
      RECT  175.3 296.0 176.3 296.8 ;
      RECT  172.9 291.6 173.9 292.4 ;
      RECT  177.3 296.0 178.1 297.6 ;
      RECT  170.5 296.0 171.3 297.6 ;
      RECT  175.1 292.8 176.3 293.6 ;
      RECT  175.5 292.4 176.3 292.8 ;
      RECT  175.5 291.6 176.5 292.4 ;
      RECT  172.9 288.4 173.7 289.2 ;
      RECT  175.7 288.4 176.5 289.2 ;
      RECT  173.1 296.0 174.1 296.8 ;
      RECT  170.5 291.2 171.3 295.4 ;
      RECT  173.1 292.4 173.9 294.6 ;
      RECT  170.5 298.4 178.1 297.6 ;
      RECT  173.1 301.4 174.7 300.6 ;
      RECT  175.5 302.4 176.3 300.0 ;
      RECT  177.3 304.8 178.1 300.6 ;
      RECT  170.5 306.2 178.1 305.4 ;
      RECT  174.3 305.4 175.1 305.2 ;
      RECT  173.1 300.6 173.9 300.0 ;
      RECT  175.3 300.0 176.3 299.2 ;
      RECT  172.9 304.4 173.9 303.6 ;
      RECT  177.3 300.0 178.1 298.4 ;
      RECT  170.5 300.0 171.3 298.4 ;
      RECT  175.1 303.2 176.3 302.4 ;
      RECT  175.5 303.6 176.3 303.2 ;
      RECT  175.5 304.4 176.5 303.6 ;
      RECT  172.9 307.6 173.7 306.8 ;
      RECT  175.7 307.6 176.5 306.8 ;
      RECT  173.1 300.0 174.1 299.2 ;
      RECT  170.5 304.8 171.3 300.6 ;
      RECT  173.1 303.6 173.9 301.4 ;
      RECT  170.5 318.4 178.1 319.2 ;
      RECT  173.1 315.4 174.7 316.2 ;
      RECT  175.5 314.4 176.3 316.8 ;
      RECT  177.3 312.0 178.1 316.2 ;
      RECT  170.5 310.6 178.1 311.4 ;
      RECT  174.3 311.4 175.1 311.6 ;
      RECT  173.1 316.2 173.9 316.8 ;
      RECT  175.3 316.8 176.3 317.6 ;
      RECT  172.9 312.4 173.9 313.2 ;
      RECT  177.3 316.8 178.1 318.4 ;
      RECT  170.5 316.8 171.3 318.4 ;
      RECT  175.1 313.6 176.3 314.4 ;
      RECT  175.5 313.2 176.3 313.6 ;
      RECT  175.5 312.4 176.5 313.2 ;
      RECT  172.9 309.2 173.7 310.0 ;
      RECT  175.7 309.2 176.5 310.0 ;
      RECT  173.1 316.8 174.1 317.6 ;
      RECT  170.5 312.0 171.3 316.2 ;
      RECT  173.1 313.2 173.9 315.4 ;
      RECT  170.5 319.2 178.1 318.4 ;
      RECT  173.1 322.2 174.7 321.4 ;
      RECT  175.5 323.2 176.3 320.8 ;
      RECT  177.3 325.6 178.1 321.4 ;
      RECT  170.5 327.0 178.1 326.2 ;
      RECT  174.3 326.2 175.1 326.0 ;
      RECT  173.1 321.4 173.9 320.8 ;
      RECT  175.3 320.8 176.3 320.0 ;
      RECT  172.9 325.2 173.9 324.4 ;
      RECT  177.3 320.8 178.1 319.2 ;
      RECT  170.5 320.8 171.3 319.2 ;
      RECT  175.1 324.0 176.3 323.2 ;
      RECT  175.5 324.4 176.3 324.0 ;
      RECT  175.5 325.2 176.5 324.4 ;
      RECT  172.9 328.4 173.7 327.6 ;
      RECT  175.7 328.4 176.5 327.6 ;
      RECT  173.1 320.8 174.1 320.0 ;
      RECT  170.5 325.6 171.3 321.4 ;
      RECT  173.1 324.4 173.9 322.2 ;
      RECT  170.5 339.2 178.1 340.0 ;
      RECT  173.1 336.2 174.7 337.0 ;
      RECT  175.5 335.2 176.3 337.6 ;
      RECT  177.3 332.8 178.1 337.0 ;
      RECT  170.5 331.4 178.1 332.2 ;
      RECT  174.3 332.2 175.1 332.4 ;
      RECT  173.1 337.0 173.9 337.6 ;
      RECT  175.3 337.6 176.3 338.4 ;
      RECT  172.9 333.2 173.9 334.0 ;
      RECT  177.3 337.6 178.1 339.2 ;
      RECT  170.5 337.6 171.3 339.2 ;
      RECT  175.1 334.4 176.3 335.2 ;
      RECT  175.5 334.0 176.3 334.4 ;
      RECT  175.5 333.2 176.5 334.0 ;
      RECT  172.9 330.0 173.7 330.8 ;
      RECT  175.7 330.0 176.5 330.8 ;
      RECT  173.1 337.6 174.1 338.4 ;
      RECT  170.5 332.8 171.3 337.0 ;
      RECT  173.1 334.0 173.9 336.2 ;
      RECT  170.5 340.0 178.1 339.2 ;
      RECT  173.1 343.0 174.7 342.2 ;
      RECT  175.5 344.0 176.3 341.6 ;
      RECT  177.3 346.4 178.1 342.2 ;
      RECT  170.5 347.8 178.1 347.0 ;
      RECT  174.3 347.0 175.1 346.8 ;
      RECT  173.1 342.2 173.9 341.6 ;
      RECT  175.3 341.6 176.3 340.8 ;
      RECT  172.9 346.0 173.9 345.2 ;
      RECT  177.3 341.6 178.1 340.0 ;
      RECT  170.5 341.6 171.3 340.0 ;
      RECT  175.1 344.8 176.3 344.0 ;
      RECT  175.5 345.2 176.3 344.8 ;
      RECT  175.5 346.0 176.5 345.2 ;
      RECT  172.9 349.2 173.7 348.4 ;
      RECT  175.7 349.2 176.5 348.4 ;
      RECT  173.1 341.6 174.1 340.8 ;
      RECT  170.5 346.4 171.3 342.2 ;
      RECT  173.1 345.2 173.9 343.0 ;
      RECT  170.5 360.0 178.1 360.8 ;
      RECT  173.1 357.0 174.7 357.8 ;
      RECT  175.5 356.0 176.3 358.4 ;
      RECT  177.3 353.6 178.1 357.8 ;
      RECT  170.5 352.2 178.1 353.0 ;
      RECT  174.3 353.0 175.1 353.2 ;
      RECT  173.1 357.8 173.9 358.4 ;
      RECT  175.3 358.4 176.3 359.2 ;
      RECT  172.9 354.0 173.9 354.8 ;
      RECT  177.3 358.4 178.1 360.0 ;
      RECT  170.5 358.4 171.3 360.0 ;
      RECT  175.1 355.2 176.3 356.0 ;
      RECT  175.5 354.8 176.3 355.2 ;
      RECT  175.5 354.0 176.5 354.8 ;
      RECT  172.9 350.8 173.7 351.6 ;
      RECT  175.7 350.8 176.5 351.6 ;
      RECT  173.1 358.4 174.1 359.2 ;
      RECT  170.5 353.6 171.3 357.8 ;
      RECT  173.1 354.8 173.9 357.0 ;
      RECT  170.9 165.0 177.7 165.8 ;
      RECT  170.9 180.6 177.7 181.4 ;
      RECT  170.9 185.8 177.7 186.6 ;
      RECT  170.9 201.4 177.7 202.2 ;
      RECT  170.9 206.6 177.7 207.4 ;
      RECT  170.9 222.2 177.7 223.0 ;
      RECT  170.9 227.4 177.7 228.2 ;
      RECT  170.9 243.0 177.7 243.8 ;
      RECT  170.9 248.2 177.7 249.0 ;
      RECT  170.9 263.8 177.7 264.6 ;
      RECT  170.9 269.0 177.7 269.8 ;
      RECT  170.9 284.6 177.7 285.4 ;
      RECT  170.9 289.8 177.7 290.6 ;
      RECT  170.9 305.4 177.7 306.2 ;
      RECT  170.9 310.6 177.7 311.4 ;
      RECT  170.9 326.2 177.7 327.0 ;
      RECT  170.9 331.4 177.7 332.2 ;
      RECT  170.9 347.0 177.7 347.8 ;
      RECT  170.9 352.2 177.7 353.0 ;
      RECT  197.7 172.8 205.3 173.6 ;
      RECT  200.3 169.8 201.9 170.6 ;
      RECT  202.7 168.8 203.5 171.2 ;
      RECT  204.5 166.4 205.3 170.6 ;
      RECT  197.7 165.0 205.3 165.8 ;
      RECT  201.5 165.8 202.3 166.0 ;
      RECT  200.3 170.6 201.1 171.2 ;
      RECT  202.5 171.2 203.5 172.0 ;
      RECT  200.1 166.8 201.1 167.6 ;
      RECT  204.5 171.2 205.3 172.8 ;
      RECT  197.7 171.2 198.5 172.8 ;
      RECT  202.3 168.0 203.5 168.8 ;
      RECT  202.7 167.6 203.5 168.0 ;
      RECT  202.7 166.8 203.7 167.6 ;
      RECT  200.1 163.6 200.9 164.4 ;
      RECT  202.9 163.6 203.7 164.4 ;
      RECT  200.3 171.2 201.3 172.0 ;
      RECT  197.7 166.4 198.5 170.6 ;
      RECT  200.3 167.6 201.1 169.8 ;
      RECT  197.7 173.6 205.3 172.8 ;
      RECT  200.3 176.6 201.9 175.8 ;
      RECT  202.7 177.6 203.5 175.2 ;
      RECT  204.5 180.0 205.3 175.8 ;
      RECT  197.7 181.4 205.3 180.6 ;
      RECT  201.5 180.6 202.3 180.4 ;
      RECT  200.3 175.8 201.1 175.2 ;
      RECT  202.5 175.2 203.5 174.4 ;
      RECT  200.1 179.6 201.1 178.8 ;
      RECT  204.5 175.2 205.3 173.6 ;
      RECT  197.7 175.2 198.5 173.6 ;
      RECT  202.3 178.4 203.5 177.6 ;
      RECT  202.7 178.8 203.5 178.4 ;
      RECT  202.7 179.6 203.7 178.8 ;
      RECT  200.1 182.8 200.9 182.0 ;
      RECT  202.9 182.8 203.7 182.0 ;
      RECT  200.3 175.2 201.3 174.4 ;
      RECT  197.7 180.0 198.5 175.8 ;
      RECT  200.3 178.8 201.1 176.6 ;
      RECT  197.7 193.6 205.3 194.4 ;
      RECT  200.3 190.6 201.9 191.4 ;
      RECT  202.7 189.6 203.5 192.0 ;
      RECT  204.5 187.2 205.3 191.4 ;
      RECT  197.7 185.8 205.3 186.6 ;
      RECT  201.5 186.6 202.3 186.8 ;
      RECT  200.3 191.4 201.1 192.0 ;
      RECT  202.5 192.0 203.5 192.8 ;
      RECT  200.1 187.6 201.1 188.4 ;
      RECT  204.5 192.0 205.3 193.6 ;
      RECT  197.7 192.0 198.5 193.6 ;
      RECT  202.3 188.8 203.5 189.6 ;
      RECT  202.7 188.4 203.5 188.8 ;
      RECT  202.7 187.6 203.7 188.4 ;
      RECT  200.1 184.4 200.9 185.2 ;
      RECT  202.9 184.4 203.7 185.2 ;
      RECT  200.3 192.0 201.3 192.8 ;
      RECT  197.7 187.2 198.5 191.4 ;
      RECT  200.3 188.4 201.1 190.6 ;
      RECT  197.7 194.4 205.3 193.6 ;
      RECT  200.3 197.4 201.9 196.6 ;
      RECT  202.7 198.4 203.5 196.0 ;
      RECT  204.5 200.8 205.3 196.6 ;
      RECT  197.7 202.2 205.3 201.4 ;
      RECT  201.5 201.4 202.3 201.2 ;
      RECT  200.3 196.6 201.1 196.0 ;
      RECT  202.5 196.0 203.5 195.2 ;
      RECT  200.1 200.4 201.1 199.6 ;
      RECT  204.5 196.0 205.3 194.4 ;
      RECT  197.7 196.0 198.5 194.4 ;
      RECT  202.3 199.2 203.5 198.4 ;
      RECT  202.7 199.6 203.5 199.2 ;
      RECT  202.7 200.4 203.7 199.6 ;
      RECT  200.1 203.6 200.9 202.8 ;
      RECT  202.9 203.6 203.7 202.8 ;
      RECT  200.3 196.0 201.3 195.2 ;
      RECT  197.7 200.8 198.5 196.6 ;
      RECT  200.3 199.6 201.1 197.4 ;
      RECT  197.7 214.4 205.3 215.2 ;
      RECT  200.3 211.4 201.9 212.2 ;
      RECT  202.7 210.4 203.5 212.8 ;
      RECT  204.5 208.0 205.3 212.2 ;
      RECT  197.7 206.6 205.3 207.4 ;
      RECT  201.5 207.4 202.3 207.6 ;
      RECT  200.3 212.2 201.1 212.8 ;
      RECT  202.5 212.8 203.5 213.6 ;
      RECT  200.1 208.4 201.1 209.2 ;
      RECT  204.5 212.8 205.3 214.4 ;
      RECT  197.7 212.8 198.5 214.4 ;
      RECT  202.3 209.6 203.5 210.4 ;
      RECT  202.7 209.2 203.5 209.6 ;
      RECT  202.7 208.4 203.7 209.2 ;
      RECT  200.1 205.2 200.9 206.0 ;
      RECT  202.9 205.2 203.7 206.0 ;
      RECT  200.3 212.8 201.3 213.6 ;
      RECT  197.7 208.0 198.5 212.2 ;
      RECT  200.3 209.2 201.1 211.4 ;
      RECT  197.7 215.2 205.3 214.4 ;
      RECT  200.3 218.2 201.9 217.4 ;
      RECT  202.7 219.2 203.5 216.8 ;
      RECT  204.5 221.6 205.3 217.4 ;
      RECT  197.7 223.0 205.3 222.2 ;
      RECT  201.5 222.2 202.3 222.0 ;
      RECT  200.3 217.4 201.1 216.8 ;
      RECT  202.5 216.8 203.5 216.0 ;
      RECT  200.1 221.2 201.1 220.4 ;
      RECT  204.5 216.8 205.3 215.2 ;
      RECT  197.7 216.8 198.5 215.2 ;
      RECT  202.3 220.0 203.5 219.2 ;
      RECT  202.7 220.4 203.5 220.0 ;
      RECT  202.7 221.2 203.7 220.4 ;
      RECT  200.1 224.4 200.9 223.6 ;
      RECT  202.9 224.4 203.7 223.6 ;
      RECT  200.3 216.8 201.3 216.0 ;
      RECT  197.7 221.6 198.5 217.4 ;
      RECT  200.3 220.4 201.1 218.2 ;
      RECT  197.7 235.2 205.3 236.0 ;
      RECT  200.3 232.2 201.9 233.0 ;
      RECT  202.7 231.2 203.5 233.6 ;
      RECT  204.5 228.8 205.3 233.0 ;
      RECT  197.7 227.4 205.3 228.2 ;
      RECT  201.5 228.2 202.3 228.4 ;
      RECT  200.3 233.0 201.1 233.6 ;
      RECT  202.5 233.6 203.5 234.4 ;
      RECT  200.1 229.2 201.1 230.0 ;
      RECT  204.5 233.6 205.3 235.2 ;
      RECT  197.7 233.6 198.5 235.2 ;
      RECT  202.3 230.4 203.5 231.2 ;
      RECT  202.7 230.0 203.5 230.4 ;
      RECT  202.7 229.2 203.7 230.0 ;
      RECT  200.1 226.0 200.9 226.8 ;
      RECT  202.9 226.0 203.7 226.8 ;
      RECT  200.3 233.6 201.3 234.4 ;
      RECT  197.7 228.8 198.5 233.0 ;
      RECT  200.3 230.0 201.1 232.2 ;
      RECT  197.7 236.0 205.3 235.2 ;
      RECT  200.3 239.0 201.9 238.2 ;
      RECT  202.7 240.0 203.5 237.6 ;
      RECT  204.5 242.4 205.3 238.2 ;
      RECT  197.7 243.8 205.3 243.0 ;
      RECT  201.5 243.0 202.3 242.8 ;
      RECT  200.3 238.2 201.1 237.6 ;
      RECT  202.5 237.6 203.5 236.8 ;
      RECT  200.1 242.0 201.1 241.2 ;
      RECT  204.5 237.6 205.3 236.0 ;
      RECT  197.7 237.6 198.5 236.0 ;
      RECT  202.3 240.8 203.5 240.0 ;
      RECT  202.7 241.2 203.5 240.8 ;
      RECT  202.7 242.0 203.7 241.2 ;
      RECT  200.1 245.2 200.9 244.4 ;
      RECT  202.9 245.2 203.7 244.4 ;
      RECT  200.3 237.6 201.3 236.8 ;
      RECT  197.7 242.4 198.5 238.2 ;
      RECT  200.3 241.2 201.1 239.0 ;
      RECT  197.7 256.0 205.3 256.8 ;
      RECT  200.3 253.0 201.9 253.8 ;
      RECT  202.7 252.0 203.5 254.4 ;
      RECT  204.5 249.6 205.3 253.8 ;
      RECT  197.7 248.2 205.3 249.0 ;
      RECT  201.5 249.0 202.3 249.2 ;
      RECT  200.3 253.8 201.1 254.4 ;
      RECT  202.5 254.4 203.5 255.2 ;
      RECT  200.1 250.0 201.1 250.8 ;
      RECT  204.5 254.4 205.3 256.0 ;
      RECT  197.7 254.4 198.5 256.0 ;
      RECT  202.3 251.2 203.5 252.0 ;
      RECT  202.7 250.8 203.5 251.2 ;
      RECT  202.7 250.0 203.7 250.8 ;
      RECT  200.1 246.8 200.9 247.6 ;
      RECT  202.9 246.8 203.7 247.6 ;
      RECT  200.3 254.4 201.3 255.2 ;
      RECT  197.7 249.6 198.5 253.8 ;
      RECT  200.3 250.8 201.1 253.0 ;
      RECT  197.7 256.8 205.3 256.0 ;
      RECT  200.3 259.8 201.9 259.0 ;
      RECT  202.7 260.8 203.5 258.4 ;
      RECT  204.5 263.2 205.3 259.0 ;
      RECT  197.7 264.6 205.3 263.8 ;
      RECT  201.5 263.8 202.3 263.6 ;
      RECT  200.3 259.0 201.1 258.4 ;
      RECT  202.5 258.4 203.5 257.6 ;
      RECT  200.1 262.8 201.1 262.0 ;
      RECT  204.5 258.4 205.3 256.8 ;
      RECT  197.7 258.4 198.5 256.8 ;
      RECT  202.3 261.6 203.5 260.8 ;
      RECT  202.7 262.0 203.5 261.6 ;
      RECT  202.7 262.8 203.7 262.0 ;
      RECT  200.1 266.0 200.9 265.2 ;
      RECT  202.9 266.0 203.7 265.2 ;
      RECT  200.3 258.4 201.3 257.6 ;
      RECT  197.7 263.2 198.5 259.0 ;
      RECT  200.3 262.0 201.1 259.8 ;
      RECT  197.7 276.8 205.3 277.6 ;
      RECT  200.3 273.8 201.9 274.6 ;
      RECT  202.7 272.8 203.5 275.2 ;
      RECT  204.5 270.4 205.3 274.6 ;
      RECT  197.7 269.0 205.3 269.8 ;
      RECT  201.5 269.8 202.3 270.0 ;
      RECT  200.3 274.6 201.1 275.2 ;
      RECT  202.5 275.2 203.5 276.0 ;
      RECT  200.1 270.8 201.1 271.6 ;
      RECT  204.5 275.2 205.3 276.8 ;
      RECT  197.7 275.2 198.5 276.8 ;
      RECT  202.3 272.0 203.5 272.8 ;
      RECT  202.7 271.6 203.5 272.0 ;
      RECT  202.7 270.8 203.7 271.6 ;
      RECT  200.1 267.6 200.9 268.4 ;
      RECT  202.9 267.6 203.7 268.4 ;
      RECT  200.3 275.2 201.3 276.0 ;
      RECT  197.7 270.4 198.5 274.6 ;
      RECT  200.3 271.6 201.1 273.8 ;
      RECT  197.7 277.6 205.3 276.8 ;
      RECT  200.3 280.6 201.9 279.8 ;
      RECT  202.7 281.6 203.5 279.2 ;
      RECT  204.5 284.0 205.3 279.8 ;
      RECT  197.7 285.4 205.3 284.6 ;
      RECT  201.5 284.6 202.3 284.4 ;
      RECT  200.3 279.8 201.1 279.2 ;
      RECT  202.5 279.2 203.5 278.4 ;
      RECT  200.1 283.6 201.1 282.8 ;
      RECT  204.5 279.2 205.3 277.6 ;
      RECT  197.7 279.2 198.5 277.6 ;
      RECT  202.3 282.4 203.5 281.6 ;
      RECT  202.7 282.8 203.5 282.4 ;
      RECT  202.7 283.6 203.7 282.8 ;
      RECT  200.1 286.8 200.9 286.0 ;
      RECT  202.9 286.8 203.7 286.0 ;
      RECT  200.3 279.2 201.3 278.4 ;
      RECT  197.7 284.0 198.5 279.8 ;
      RECT  200.3 282.8 201.1 280.6 ;
      RECT  197.7 297.6 205.3 298.4 ;
      RECT  200.3 294.6 201.9 295.4 ;
      RECT  202.7 293.6 203.5 296.0 ;
      RECT  204.5 291.2 205.3 295.4 ;
      RECT  197.7 289.8 205.3 290.6 ;
      RECT  201.5 290.6 202.3 290.8 ;
      RECT  200.3 295.4 201.1 296.0 ;
      RECT  202.5 296.0 203.5 296.8 ;
      RECT  200.1 291.6 201.1 292.4 ;
      RECT  204.5 296.0 205.3 297.6 ;
      RECT  197.7 296.0 198.5 297.6 ;
      RECT  202.3 292.8 203.5 293.6 ;
      RECT  202.7 292.4 203.5 292.8 ;
      RECT  202.7 291.6 203.7 292.4 ;
      RECT  200.1 288.4 200.9 289.2 ;
      RECT  202.9 288.4 203.7 289.2 ;
      RECT  200.3 296.0 201.3 296.8 ;
      RECT  197.7 291.2 198.5 295.4 ;
      RECT  200.3 292.4 201.1 294.6 ;
      RECT  197.7 298.4 205.3 297.6 ;
      RECT  200.3 301.4 201.9 300.6 ;
      RECT  202.7 302.4 203.5 300.0 ;
      RECT  204.5 304.8 205.3 300.6 ;
      RECT  197.7 306.2 205.3 305.4 ;
      RECT  201.5 305.4 202.3 305.2 ;
      RECT  200.3 300.6 201.1 300.0 ;
      RECT  202.5 300.0 203.5 299.2 ;
      RECT  200.1 304.4 201.1 303.6 ;
      RECT  204.5 300.0 205.3 298.4 ;
      RECT  197.7 300.0 198.5 298.4 ;
      RECT  202.3 303.2 203.5 302.4 ;
      RECT  202.7 303.6 203.5 303.2 ;
      RECT  202.7 304.4 203.7 303.6 ;
      RECT  200.1 307.6 200.9 306.8 ;
      RECT  202.9 307.6 203.7 306.8 ;
      RECT  200.3 300.0 201.3 299.2 ;
      RECT  197.7 304.8 198.5 300.6 ;
      RECT  200.3 303.6 201.1 301.4 ;
      RECT  197.7 318.4 205.3 319.2 ;
      RECT  200.3 315.4 201.9 316.2 ;
      RECT  202.7 314.4 203.5 316.8 ;
      RECT  204.5 312.0 205.3 316.2 ;
      RECT  197.7 310.6 205.3 311.4 ;
      RECT  201.5 311.4 202.3 311.6 ;
      RECT  200.3 316.2 201.1 316.8 ;
      RECT  202.5 316.8 203.5 317.6 ;
      RECT  200.1 312.4 201.1 313.2 ;
      RECT  204.5 316.8 205.3 318.4 ;
      RECT  197.7 316.8 198.5 318.4 ;
      RECT  202.3 313.6 203.5 314.4 ;
      RECT  202.7 313.2 203.5 313.6 ;
      RECT  202.7 312.4 203.7 313.2 ;
      RECT  200.1 309.2 200.9 310.0 ;
      RECT  202.9 309.2 203.7 310.0 ;
      RECT  200.3 316.8 201.3 317.6 ;
      RECT  197.7 312.0 198.5 316.2 ;
      RECT  200.3 313.2 201.1 315.4 ;
      RECT  197.7 319.2 205.3 318.4 ;
      RECT  200.3 322.2 201.9 321.4 ;
      RECT  202.7 323.2 203.5 320.8 ;
      RECT  204.5 325.6 205.3 321.4 ;
      RECT  197.7 327.0 205.3 326.2 ;
      RECT  201.5 326.2 202.3 326.0 ;
      RECT  200.3 321.4 201.1 320.8 ;
      RECT  202.5 320.8 203.5 320.0 ;
      RECT  200.1 325.2 201.1 324.4 ;
      RECT  204.5 320.8 205.3 319.2 ;
      RECT  197.7 320.8 198.5 319.2 ;
      RECT  202.3 324.0 203.5 323.2 ;
      RECT  202.7 324.4 203.5 324.0 ;
      RECT  202.7 325.2 203.7 324.4 ;
      RECT  200.1 328.4 200.9 327.6 ;
      RECT  202.9 328.4 203.7 327.6 ;
      RECT  200.3 320.8 201.3 320.0 ;
      RECT  197.7 325.6 198.5 321.4 ;
      RECT  200.3 324.4 201.1 322.2 ;
      RECT  197.7 339.2 205.3 340.0 ;
      RECT  200.3 336.2 201.9 337.0 ;
      RECT  202.7 335.2 203.5 337.6 ;
      RECT  204.5 332.8 205.3 337.0 ;
      RECT  197.7 331.4 205.3 332.2 ;
      RECT  201.5 332.2 202.3 332.4 ;
      RECT  200.3 337.0 201.1 337.6 ;
      RECT  202.5 337.6 203.5 338.4 ;
      RECT  200.1 333.2 201.1 334.0 ;
      RECT  204.5 337.6 205.3 339.2 ;
      RECT  197.7 337.6 198.5 339.2 ;
      RECT  202.3 334.4 203.5 335.2 ;
      RECT  202.7 334.0 203.5 334.4 ;
      RECT  202.7 333.2 203.7 334.0 ;
      RECT  200.1 330.0 200.9 330.8 ;
      RECT  202.9 330.0 203.7 330.8 ;
      RECT  200.3 337.6 201.3 338.4 ;
      RECT  197.7 332.8 198.5 337.0 ;
      RECT  200.3 334.0 201.1 336.2 ;
      RECT  197.7 340.0 205.3 339.2 ;
      RECT  200.3 343.0 201.9 342.2 ;
      RECT  202.7 344.0 203.5 341.6 ;
      RECT  204.5 346.4 205.3 342.2 ;
      RECT  197.7 347.8 205.3 347.0 ;
      RECT  201.5 347.0 202.3 346.8 ;
      RECT  200.3 342.2 201.1 341.6 ;
      RECT  202.5 341.6 203.5 340.8 ;
      RECT  200.1 346.0 201.1 345.2 ;
      RECT  204.5 341.6 205.3 340.0 ;
      RECT  197.7 341.6 198.5 340.0 ;
      RECT  202.3 344.8 203.5 344.0 ;
      RECT  202.7 345.2 203.5 344.8 ;
      RECT  202.7 346.0 203.7 345.2 ;
      RECT  200.1 349.2 200.9 348.4 ;
      RECT  202.9 349.2 203.7 348.4 ;
      RECT  200.3 341.6 201.3 340.8 ;
      RECT  197.7 346.4 198.5 342.2 ;
      RECT  200.3 345.2 201.1 343.0 ;
      RECT  197.7 360.0 205.3 360.8 ;
      RECT  200.3 357.0 201.9 357.8 ;
      RECT  202.7 356.0 203.5 358.4 ;
      RECT  204.5 353.6 205.3 357.8 ;
      RECT  197.7 352.2 205.3 353.0 ;
      RECT  201.5 353.0 202.3 353.2 ;
      RECT  200.3 357.8 201.1 358.4 ;
      RECT  202.5 358.4 203.5 359.2 ;
      RECT  200.1 354.0 201.1 354.8 ;
      RECT  204.5 358.4 205.3 360.0 ;
      RECT  197.7 358.4 198.5 360.0 ;
      RECT  202.3 355.2 203.5 356.0 ;
      RECT  202.7 354.8 203.5 355.2 ;
      RECT  202.7 354.0 203.7 354.8 ;
      RECT  200.1 350.8 200.9 351.6 ;
      RECT  202.9 350.8 203.7 351.6 ;
      RECT  200.3 358.4 201.3 359.2 ;
      RECT  197.7 353.6 198.5 357.8 ;
      RECT  200.3 354.8 201.1 357.0 ;
      RECT  198.1 165.0 204.9 165.8 ;
      RECT  198.1 180.6 204.9 181.4 ;
      RECT  198.1 185.8 204.9 186.6 ;
      RECT  198.1 201.4 204.9 202.2 ;
      RECT  198.1 206.6 204.9 207.4 ;
      RECT  198.1 222.2 204.9 223.0 ;
      RECT  198.1 227.4 204.9 228.2 ;
      RECT  198.1 243.0 204.9 243.8 ;
      RECT  198.1 248.2 204.9 249.0 ;
      RECT  198.1 263.8 204.9 264.6 ;
      RECT  198.1 269.0 204.9 269.8 ;
      RECT  198.1 284.6 204.9 285.4 ;
      RECT  198.1 289.8 204.9 290.6 ;
      RECT  198.1 305.4 204.9 306.2 ;
      RECT  198.1 310.6 204.9 311.4 ;
      RECT  198.1 326.2 204.9 327.0 ;
      RECT  198.1 331.4 204.9 332.2 ;
      RECT  198.1 347.0 204.9 347.8 ;
      RECT  198.1 352.2 204.9 353.0 ;
      RECT  170.9 185.8 204.9 186.6 ;
      RECT  170.9 201.4 204.9 202.2 ;
      RECT  170.9 206.6 204.9 207.4 ;
      RECT  170.9 222.2 204.9 223.0 ;
      RECT  170.9 227.4 204.9 228.2 ;
      RECT  170.9 243.0 204.9 243.8 ;
      RECT  170.9 248.2 204.9 249.0 ;
      RECT  170.9 263.8 204.9 264.6 ;
      RECT  170.9 269.0 204.9 269.8 ;
      RECT  170.9 284.6 204.9 285.4 ;
      RECT  170.9 289.8 204.9 290.6 ;
      RECT  170.9 305.4 204.9 306.2 ;
      RECT  170.9 310.6 204.9 311.4 ;
      RECT  170.9 326.2 204.9 327.0 ;
      RECT  170.9 331.4 204.9 332.2 ;
      RECT  170.9 347.0 204.9 347.8 ;
      RECT  170.9 180.6 204.9 181.4 ;
      RECT  181.2 149.6 182.0 150.4 ;
      RECT  179.2 149.6 180.0 150.4 ;
      RECT  181.2 154.0 182.0 154.8 ;
      RECT  179.2 154.0 180.0 154.8 ;
      RECT  183.2 154.0 184.0 154.8 ;
      RECT  181.2 154.0 182.0 154.8 ;
      RECT  177.7 147.5 184.5 148.1 ;
      RECT  188.0 149.6 188.8 150.4 ;
      RECT  186.0 149.6 186.8 150.4 ;
      RECT  188.0 154.0 188.8 154.8 ;
      RECT  186.0 154.0 186.8 154.8 ;
      RECT  190.0 154.0 190.8 154.8 ;
      RECT  188.0 154.0 188.8 154.8 ;
      RECT  184.5 147.5 191.3 148.1 ;
      RECT  194.8 149.6 195.6 150.4 ;
      RECT  192.8 149.6 193.6 150.4 ;
      RECT  194.8 154.0 195.6 154.8 ;
      RECT  192.8 154.0 193.6 154.8 ;
      RECT  196.8 154.0 197.6 154.8 ;
      RECT  194.8 154.0 195.6 154.8 ;
      RECT  191.3 147.5 198.1 148.1 ;
      RECT  177.7 147.5 198.1 148.1 ;
      RECT  189.1 130.8 189.9 133.2 ;
      RECT  185.7 120.0 187.1 120.6 ;
      RECT  187.5 131.4 188.3 133.2 ;
      RECT  189.9 123.0 190.7 124.2 ;
      RECT  185.7 118.6 186.3 120.0 ;
      RECT  185.1 113.8 186.5 114.4 ;
      RECT  190.7 118.6 191.3 120.0 ;
      RECT  187.7 135.8 188.5 137.6 ;
      RECT  184.1 139.6 191.7 140.4 ;
      RECT  186.3 120.6 187.1 120.8 ;
      RECT  185.7 114.4 186.5 118.6 ;
      RECT  185.9 122.8 187.1 123.6 ;
      RECT  188.9 113.8 189.7 119.4 ;
      RECT  187.5 124.2 190.7 124.8 ;
      RECT  187.1 118.6 187.9 119.4 ;
      RECT  189.1 130.0 190.5 130.8 ;
      RECT  190.9 137.2 191.7 138.0 ;
      RECT  189.3 136.4 191.7 137.2 ;
      RECT  187.7 133.2 188.3 135.8 ;
      RECT  187.3 113.8 188.1 118.6 ;
      RECT  190.5 113.8 191.3 118.6 ;
      RECT  190.3 120.0 191.3 120.8 ;
      RECT  189.1 125.4 189.9 130.0 ;
      RECT  185.1 112.0 185.9 113.8 ;
      RECT  189.3 137.2 190.1 137.6 ;
      RECT  185.9 123.6 186.7 133.2 ;
      RECT  187.5 124.8 188.1 125.4 ;
      RECT  189.3 135.8 190.1 136.4 ;
      RECT  187.5 125.4 188.3 129.0 ;
      RECT  195.9 130.8 196.7 133.2 ;
      RECT  192.5 120.0 193.9 120.6 ;
      RECT  194.3 131.4 195.1 133.2 ;
      RECT  196.7 123.0 197.5 124.2 ;
      RECT  192.5 118.6 193.1 120.0 ;
      RECT  191.9 113.8 193.3 114.4 ;
      RECT  197.5 118.6 198.1 120.0 ;
      RECT  194.5 135.8 195.3 137.6 ;
      RECT  190.9 139.6 198.5 140.4 ;
      RECT  193.1 120.6 193.9 120.8 ;
      RECT  192.5 114.4 193.3 118.6 ;
      RECT  192.7 122.8 193.9 123.6 ;
      RECT  195.7 113.8 196.5 119.4 ;
      RECT  194.3 124.2 197.5 124.8 ;
      RECT  193.9 118.6 194.7 119.4 ;
      RECT  195.9 130.0 197.3 130.8 ;
      RECT  197.7 137.2 198.5 138.0 ;
      RECT  196.1 136.4 198.5 137.2 ;
      RECT  194.5 133.2 195.1 135.8 ;
      RECT  194.1 113.8 194.9 118.6 ;
      RECT  197.3 113.8 198.1 118.6 ;
      RECT  197.1 120.0 198.1 120.8 ;
      RECT  195.9 125.4 196.7 130.0 ;
      RECT  191.9 112.0 192.7 113.8 ;
      RECT  196.1 137.2 196.9 137.6 ;
      RECT  192.7 123.6 193.5 133.2 ;
      RECT  194.3 124.8 194.9 125.4 ;
      RECT  196.1 135.8 196.9 136.4 ;
      RECT  194.3 125.4 195.1 129.0 ;
      RECT  184.5 139.7 198.1 140.3 ;
      RECT  188.3 76.4 189.1 78.6 ;
      RECT  186.9 88.6 188.5 89.4 ;
      RECT  188.7 84.2 189.9 85.0 ;
      RECT  185.5 81.4 186.3 85.2 ;
      RECT  186.9 89.4 187.7 91.4 ;
      RECT  188.7 81.4 190.5 82.8 ;
      RECT  189.1 80.0 190.7 80.8 ;
      RECT  185.5 85.2 189.5 85.8 ;
      RECT  188.7 85.0 189.5 85.2 ;
      RECT  186.7 76.4 187.5 77.8 ;
      RECT  185.3 100.6 186.1 103.0 ;
      RECT  185.5 85.8 186.3 87.8 ;
      RECT  188.7 85.8 189.5 87.8 ;
      RECT  186.7 72.6 187.5 74.6 ;
      RECT  187.1 81.4 187.9 82.8 ;
      RECT  185.1 75.2 185.9 77.8 ;
      RECT  188.5 93.4 189.3 94.6 ;
      RECT  185.1 79.2 185.9 80.0 ;
      RECT  185.1 71.2 189.1 72.0 ;
      RECT  187.5 66.2 188.3 67.8 ;
      RECT  188.5 90.0 189.3 92.6 ;
      RECT  188.5 100.6 189.3 103.8 ;
      RECT  185.1 72.0 185.9 74.0 ;
      RECT  188.3 72.0 189.1 74.0 ;
      RECT  188.5 92.6 191.1 93.4 ;
      RECT  190.1 101.4 191.1 102.2 ;
      RECT  185.3 90.0 186.1 98.6 ;
      RECT  185.1 74.6 187.5 75.2 ;
      RECT  186.9 93.8 187.7 103.0 ;
      RECT  189.5 82.8 190.5 83.0 ;
      RECT  185.1 69.8 190.7 70.6 ;
      RECT  190.5 93.4 191.1 101.4 ;
      RECT  187.1 86.4 187.9 88.6 ;
      RECT  189.9 72.6 190.7 80.0 ;
      RECT  185.5 103.0 186.1 103.6 ;
      RECT  185.3 77.8 185.9 79.2 ;
      RECT  185.5 103.6 187.3 104.4 ;
      RECT  195.1 76.4 195.9 78.6 ;
      RECT  193.7 88.6 195.3 89.4 ;
      RECT  195.5 84.2 196.7 85.0 ;
      RECT  192.3 81.4 193.1 85.2 ;
      RECT  193.7 89.4 194.5 91.4 ;
      RECT  195.5 81.4 197.3 82.8 ;
      RECT  195.9 80.0 197.5 80.8 ;
      RECT  192.3 85.2 196.3 85.8 ;
      RECT  195.5 85.0 196.3 85.2 ;
      RECT  193.5 76.4 194.3 77.8 ;
      RECT  192.1 100.6 192.9 103.0 ;
      RECT  192.3 85.8 193.1 87.8 ;
      RECT  195.5 85.8 196.3 87.8 ;
      RECT  193.5 72.6 194.3 74.6 ;
      RECT  193.9 81.4 194.7 82.8 ;
      RECT  191.9 75.2 192.7 77.8 ;
      RECT  195.3 93.4 196.1 94.6 ;
      RECT  191.9 79.2 192.7 80.0 ;
      RECT  191.9 71.2 195.9 72.0 ;
      RECT  194.3 66.2 195.1 67.8 ;
      RECT  195.3 90.0 196.1 92.6 ;
      RECT  195.3 100.6 196.1 103.8 ;
      RECT  191.9 72.0 192.7 74.0 ;
      RECT  195.1 72.0 195.9 74.0 ;
      RECT  195.3 92.6 197.9 93.4 ;
      RECT  196.9 101.4 197.9 102.2 ;
      RECT  192.1 90.0 192.9 98.6 ;
      RECT  191.9 74.6 194.3 75.2 ;
      RECT  193.7 93.8 194.5 103.0 ;
      RECT  196.3 82.8 197.3 83.0 ;
      RECT  191.9 69.8 197.5 70.6 ;
      RECT  197.3 93.4 197.9 101.4 ;
      RECT  193.9 86.4 194.7 88.6 ;
      RECT  196.7 72.6 197.5 80.0 ;
      RECT  192.3 103.0 192.9 103.6 ;
      RECT  192.1 77.8 192.7 79.2 ;
      RECT  192.3 103.6 194.1 104.4 ;
      RECT  184.5 69.8 198.1 70.4 ;
      RECT  184.5 140.3 198.1 139.7 ;
      RECT  177.7 148.1 198.1 147.5 ;
      RECT  184.5 70.4 198.1 69.8 ;
      RECT  94.9 192.3 95.7 193.1 ;
      RECT  92.9 192.3 93.7 193.1 ;
      RECT  94.9 184.9 95.7 185.7 ;
      RECT  92.9 184.9 93.7 185.7 ;
      RECT  93.3 188.6 94.1 189.4 ;
      RECT  95.3 188.7 95.9 189.3 ;
      RECT  91.7 194.1 98.3 194.7 ;
      RECT  91.7 183.7 98.3 184.3 ;
      RECT  94.9 196.5 95.7 195.7 ;
      RECT  92.9 196.5 93.7 195.7 ;
      RECT  94.9 203.9 95.7 203.1 ;
      RECT  92.9 203.9 93.7 203.1 ;
      RECT  93.3 200.2 94.1 199.4 ;
      RECT  95.3 200.1 95.9 199.5 ;
      RECT  91.7 194.7 98.3 194.1 ;
      RECT  91.7 205.1 98.3 204.5 ;
      RECT  109.9 192.3 110.7 193.1 ;
      RECT  107.9 192.3 108.7 193.1 ;
      RECT  111.9 192.3 112.7 193.1 ;
      RECT  109.9 192.3 110.7 193.1 ;
      RECT  107.9 185.3 108.7 186.1 ;
      RECT  111.9 185.3 112.7 186.1 ;
      RECT  108.9 186.8 109.7 187.6 ;
      RECT  110.9 189.6 111.7 190.4 ;
      RECT  113.4 191.0 114.0 191.6 ;
      RECT  106.7 194.1 115.3 194.7 ;
      RECT  106.7 183.7 115.3 184.3 ;
      RECT  118.5 192.3 119.3 193.1 ;
      RECT  116.5 192.3 117.3 193.1 ;
      RECT  118.5 184.9 119.3 185.7 ;
      RECT  116.5 184.9 117.3 185.7 ;
      RECT  116.9 188.6 117.7 189.4 ;
      RECT  118.9 188.7 119.5 189.3 ;
      RECT  115.3 194.1 121.9 194.7 ;
      RECT  115.3 183.7 121.9 184.3 ;
      RECT  108.9 186.8 109.7 187.6 ;
      RECT  110.9 189.6 111.7 190.4 ;
      RECT  118.9 188.7 119.5 189.3 ;
      RECT  106.7 194.1 121.9 194.7 ;
      RECT  106.7 183.7 121.9 184.3 ;
      RECT  109.9 196.5 110.7 195.7 ;
      RECT  107.9 196.5 108.7 195.7 ;
      RECT  111.9 196.5 112.7 195.7 ;
      RECT  109.9 196.5 110.7 195.7 ;
      RECT  107.9 203.5 108.7 202.7 ;
      RECT  111.9 203.5 112.7 202.7 ;
      RECT  108.9 202.0 109.7 201.2 ;
      RECT  110.9 199.2 111.7 198.4 ;
      RECT  113.4 197.8 114.0 197.2 ;
      RECT  106.7 194.7 115.3 194.1 ;
      RECT  106.7 205.1 115.3 204.5 ;
      RECT  118.5 196.5 119.3 195.7 ;
      RECT  116.5 196.5 117.3 195.7 ;
      RECT  118.5 203.9 119.3 203.1 ;
      RECT  116.5 203.9 117.3 203.1 ;
      RECT  116.9 200.2 117.7 199.4 ;
      RECT  118.9 200.1 119.5 199.5 ;
      RECT  115.3 194.7 121.9 194.1 ;
      RECT  115.3 205.1 121.9 204.5 ;
      RECT  108.9 202.0 109.7 201.2 ;
      RECT  110.9 199.2 111.7 198.4 ;
      RECT  118.9 200.1 119.5 199.5 ;
      RECT  106.7 194.7 121.9 194.1 ;
      RECT  106.7 205.1 121.9 204.5 ;
      RECT  109.9 213.1 110.7 213.9 ;
      RECT  107.9 213.1 108.7 213.9 ;
      RECT  111.9 213.1 112.7 213.9 ;
      RECT  109.9 213.1 110.7 213.9 ;
      RECT  107.9 206.1 108.7 206.9 ;
      RECT  111.9 206.1 112.7 206.9 ;
      RECT  108.9 207.6 109.7 208.4 ;
      RECT  110.9 210.4 111.7 211.2 ;
      RECT  113.4 211.8 114.0 212.4 ;
      RECT  106.7 214.9 115.3 215.5 ;
      RECT  106.7 204.5 115.3 205.1 ;
      RECT  118.5 213.1 119.3 213.9 ;
      RECT  116.5 213.1 117.3 213.9 ;
      RECT  118.5 205.7 119.3 206.5 ;
      RECT  116.5 205.7 117.3 206.5 ;
      RECT  116.9 209.4 117.7 210.2 ;
      RECT  118.9 209.5 119.5 210.1 ;
      RECT  115.3 214.9 121.9 215.5 ;
      RECT  115.3 204.5 121.9 205.1 ;
      RECT  108.9 207.6 109.7 208.4 ;
      RECT  110.9 210.4 111.7 211.2 ;
      RECT  118.9 209.5 119.5 210.1 ;
      RECT  106.7 214.9 121.9 215.5 ;
      RECT  106.7 204.5 121.9 205.1 ;
      RECT  109.9 217.3 110.7 216.5 ;
      RECT  107.9 217.3 108.7 216.5 ;
      RECT  111.9 217.3 112.7 216.5 ;
      RECT  109.9 217.3 110.7 216.5 ;
      RECT  107.9 224.3 108.7 223.5 ;
      RECT  111.9 224.3 112.7 223.5 ;
      RECT  108.9 222.8 109.7 222.0 ;
      RECT  110.9 220.0 111.7 219.2 ;
      RECT  113.4 218.6 114.0 218.0 ;
      RECT  106.7 215.5 115.3 214.9 ;
      RECT  106.7 225.9 115.3 225.3 ;
      RECT  118.5 217.3 119.3 216.5 ;
      RECT  116.5 217.3 117.3 216.5 ;
      RECT  118.5 224.7 119.3 223.9 ;
      RECT  116.5 224.7 117.3 223.9 ;
      RECT  116.9 221.0 117.7 220.2 ;
      RECT  118.9 220.9 119.5 220.3 ;
      RECT  115.3 215.5 121.9 214.9 ;
      RECT  115.3 225.9 121.9 225.3 ;
      RECT  108.9 222.8 109.7 222.0 ;
      RECT  110.9 220.0 111.7 219.2 ;
      RECT  118.9 220.9 119.5 220.3 ;
      RECT  106.7 215.5 121.9 214.9 ;
      RECT  106.7 225.9 121.9 225.3 ;
      RECT  118.9 188.7 119.5 189.3 ;
      RECT  118.9 199.5 119.5 200.1 ;
      RECT  118.9 209.5 119.5 210.1 ;
      RECT  118.9 220.3 119.5 220.9 ;
      RECT  94.9 254.7 95.7 255.5 ;
      RECT  92.9 254.7 93.7 255.5 ;
      RECT  94.9 247.3 95.7 248.1 ;
      RECT  92.9 247.3 93.7 248.1 ;
      RECT  93.3 251.0 94.1 251.8 ;
      RECT  95.3 251.1 95.9 251.7 ;
      RECT  91.7 256.5 98.3 257.1 ;
      RECT  91.7 246.1 98.3 246.7 ;
      RECT  94.9 258.9 95.7 258.1 ;
      RECT  92.9 258.9 93.7 258.1 ;
      RECT  94.9 266.3 95.7 265.5 ;
      RECT  92.9 266.3 93.7 265.5 ;
      RECT  93.3 262.6 94.1 261.8 ;
      RECT  95.3 262.5 95.9 261.9 ;
      RECT  91.7 257.1 98.3 256.5 ;
      RECT  91.7 267.5 98.3 266.9 ;
      RECT  109.9 254.7 110.7 255.5 ;
      RECT  107.9 254.7 108.7 255.5 ;
      RECT  111.9 254.7 112.7 255.5 ;
      RECT  109.9 254.7 110.7 255.5 ;
      RECT  107.9 247.7 108.7 248.5 ;
      RECT  111.9 247.7 112.7 248.5 ;
      RECT  108.9 249.2 109.7 250.0 ;
      RECT  110.9 252.0 111.7 252.8 ;
      RECT  113.4 253.4 114.0 254.0 ;
      RECT  106.7 256.5 115.3 257.1 ;
      RECT  106.7 246.1 115.3 246.7 ;
      RECT  118.5 254.7 119.3 255.5 ;
      RECT  116.5 254.7 117.3 255.5 ;
      RECT  118.5 247.3 119.3 248.1 ;
      RECT  116.5 247.3 117.3 248.1 ;
      RECT  116.9 251.0 117.7 251.8 ;
      RECT  118.9 251.1 119.5 251.7 ;
      RECT  115.3 256.5 121.9 257.1 ;
      RECT  115.3 246.1 121.9 246.7 ;
      RECT  108.9 249.2 109.7 250.0 ;
      RECT  110.9 252.0 111.7 252.8 ;
      RECT  118.9 251.1 119.5 251.7 ;
      RECT  106.7 256.5 121.9 257.1 ;
      RECT  106.7 246.1 121.9 246.7 ;
      RECT  109.9 258.9 110.7 258.1 ;
      RECT  107.9 258.9 108.7 258.1 ;
      RECT  111.9 258.9 112.7 258.1 ;
      RECT  109.9 258.9 110.7 258.1 ;
      RECT  107.9 265.9 108.7 265.1 ;
      RECT  111.9 265.9 112.7 265.1 ;
      RECT  108.9 264.4 109.7 263.6 ;
      RECT  110.9 261.6 111.7 260.8 ;
      RECT  113.4 260.2 114.0 259.6 ;
      RECT  106.7 257.1 115.3 256.5 ;
      RECT  106.7 267.5 115.3 266.9 ;
      RECT  118.5 258.9 119.3 258.1 ;
      RECT  116.5 258.9 117.3 258.1 ;
      RECT  118.5 266.3 119.3 265.5 ;
      RECT  116.5 266.3 117.3 265.5 ;
      RECT  116.9 262.6 117.7 261.8 ;
      RECT  118.9 262.5 119.5 261.9 ;
      RECT  115.3 257.1 121.9 256.5 ;
      RECT  115.3 267.5 121.9 266.9 ;
      RECT  108.9 264.4 109.7 263.6 ;
      RECT  110.9 261.6 111.7 260.8 ;
      RECT  118.9 262.5 119.5 261.9 ;
      RECT  106.7 257.1 121.9 256.5 ;
      RECT  106.7 267.5 121.9 266.9 ;
      RECT  109.9 275.5 110.7 276.3 ;
      RECT  107.9 275.5 108.7 276.3 ;
      RECT  111.9 275.5 112.7 276.3 ;
      RECT  109.9 275.5 110.7 276.3 ;
      RECT  107.9 268.5 108.7 269.3 ;
      RECT  111.9 268.5 112.7 269.3 ;
      RECT  108.9 270.0 109.7 270.8 ;
      RECT  110.9 272.8 111.7 273.6 ;
      RECT  113.4 274.2 114.0 274.8 ;
      RECT  106.7 277.3 115.3 277.9 ;
      RECT  106.7 266.9 115.3 267.5 ;
      RECT  118.5 275.5 119.3 276.3 ;
      RECT  116.5 275.5 117.3 276.3 ;
      RECT  118.5 268.1 119.3 268.9 ;
      RECT  116.5 268.1 117.3 268.9 ;
      RECT  116.9 271.8 117.7 272.6 ;
      RECT  118.9 271.9 119.5 272.5 ;
      RECT  115.3 277.3 121.9 277.9 ;
      RECT  115.3 266.9 121.9 267.5 ;
      RECT  108.9 270.0 109.7 270.8 ;
      RECT  110.9 272.8 111.7 273.6 ;
      RECT  118.9 271.9 119.5 272.5 ;
      RECT  106.7 277.3 121.9 277.9 ;
      RECT  106.7 266.9 121.9 267.5 ;
      RECT  109.9 279.7 110.7 278.9 ;
      RECT  107.9 279.7 108.7 278.9 ;
      RECT  111.9 279.7 112.7 278.9 ;
      RECT  109.9 279.7 110.7 278.9 ;
      RECT  107.9 286.7 108.7 285.9 ;
      RECT  111.9 286.7 112.7 285.9 ;
      RECT  108.9 285.2 109.7 284.4 ;
      RECT  110.9 282.4 111.7 281.6 ;
      RECT  113.4 281.0 114.0 280.4 ;
      RECT  106.7 277.9 115.3 277.3 ;
      RECT  106.7 288.3 115.3 287.7 ;
      RECT  118.5 279.7 119.3 278.9 ;
      RECT  116.5 279.7 117.3 278.9 ;
      RECT  118.5 287.1 119.3 286.3 ;
      RECT  116.5 287.1 117.3 286.3 ;
      RECT  116.9 283.4 117.7 282.6 ;
      RECT  118.9 283.3 119.5 282.7 ;
      RECT  115.3 277.9 121.9 277.3 ;
      RECT  115.3 288.3 121.9 287.7 ;
      RECT  108.9 285.2 109.7 284.4 ;
      RECT  110.9 282.4 111.7 281.6 ;
      RECT  118.9 283.3 119.5 282.7 ;
      RECT  106.7 277.9 121.9 277.3 ;
      RECT  106.7 288.3 121.9 287.7 ;
      RECT  118.9 251.1 119.5 251.7 ;
      RECT  118.9 261.9 119.5 262.5 ;
      RECT  118.9 271.9 119.5 272.5 ;
      RECT  118.9 282.7 119.5 283.3 ;
      RECT  137.7 192.3 138.5 193.1 ;
      RECT  135.7 192.3 136.5 193.1 ;
      RECT  139.7 192.3 140.5 193.1 ;
      RECT  137.7 192.3 138.5 193.1 ;
      RECT  135.7 185.3 136.5 186.1 ;
      RECT  139.7 185.3 140.5 186.1 ;
      RECT  136.7 186.8 137.5 187.6 ;
      RECT  138.7 189.6 139.5 190.4 ;
      RECT  141.2 191.0 141.8 191.6 ;
      RECT  134.5 194.1 143.1 194.7 ;
      RECT  134.5 183.7 143.1 184.3 ;
      RECT  146.3 192.3 147.1 193.1 ;
      RECT  144.3 192.3 145.1 193.1 ;
      RECT  146.3 184.9 147.1 185.7 ;
      RECT  144.3 184.9 145.1 185.7 ;
      RECT  144.7 188.6 145.5 189.4 ;
      RECT  146.7 188.7 147.3 189.3 ;
      RECT  143.1 194.1 149.7 194.7 ;
      RECT  143.1 183.7 149.7 184.3 ;
      RECT  136.7 186.8 137.5 187.6 ;
      RECT  138.7 189.6 139.5 190.4 ;
      RECT  146.7 188.7 147.3 189.3 ;
      RECT  134.5 194.1 149.7 194.7 ;
      RECT  134.5 183.7 149.7 184.3 ;
      RECT  137.7 196.5 138.5 195.7 ;
      RECT  135.7 196.5 136.5 195.7 ;
      RECT  139.7 196.5 140.5 195.7 ;
      RECT  137.7 196.5 138.5 195.7 ;
      RECT  135.7 203.5 136.5 202.7 ;
      RECT  139.7 203.5 140.5 202.7 ;
      RECT  136.7 202.0 137.5 201.2 ;
      RECT  138.7 199.2 139.5 198.4 ;
      RECT  141.2 197.8 141.8 197.2 ;
      RECT  134.5 194.7 143.1 194.1 ;
      RECT  134.5 205.1 143.1 204.5 ;
      RECT  146.3 196.5 147.1 195.7 ;
      RECT  144.3 196.5 145.1 195.7 ;
      RECT  146.3 203.9 147.1 203.1 ;
      RECT  144.3 203.9 145.1 203.1 ;
      RECT  144.7 200.2 145.5 199.4 ;
      RECT  146.7 200.1 147.3 199.5 ;
      RECT  143.1 194.7 149.7 194.1 ;
      RECT  143.1 205.1 149.7 204.5 ;
      RECT  136.7 202.0 137.5 201.2 ;
      RECT  138.7 199.2 139.5 198.4 ;
      RECT  146.7 200.1 147.3 199.5 ;
      RECT  134.5 194.7 149.7 194.1 ;
      RECT  134.5 205.1 149.7 204.5 ;
      RECT  137.7 213.1 138.5 213.9 ;
      RECT  135.7 213.1 136.5 213.9 ;
      RECT  139.7 213.1 140.5 213.9 ;
      RECT  137.7 213.1 138.5 213.9 ;
      RECT  135.7 206.1 136.5 206.9 ;
      RECT  139.7 206.1 140.5 206.9 ;
      RECT  136.7 207.6 137.5 208.4 ;
      RECT  138.7 210.4 139.5 211.2 ;
      RECT  141.2 211.8 141.8 212.4 ;
      RECT  134.5 214.9 143.1 215.5 ;
      RECT  134.5 204.5 143.1 205.1 ;
      RECT  146.3 213.1 147.1 213.9 ;
      RECT  144.3 213.1 145.1 213.9 ;
      RECT  146.3 205.7 147.1 206.5 ;
      RECT  144.3 205.7 145.1 206.5 ;
      RECT  144.7 209.4 145.5 210.2 ;
      RECT  146.7 209.5 147.3 210.1 ;
      RECT  143.1 214.9 149.7 215.5 ;
      RECT  143.1 204.5 149.7 205.1 ;
      RECT  136.7 207.6 137.5 208.4 ;
      RECT  138.7 210.4 139.5 211.2 ;
      RECT  146.7 209.5 147.3 210.1 ;
      RECT  134.5 214.9 149.7 215.5 ;
      RECT  134.5 204.5 149.7 205.1 ;
      RECT  137.7 217.3 138.5 216.5 ;
      RECT  135.7 217.3 136.5 216.5 ;
      RECT  139.7 217.3 140.5 216.5 ;
      RECT  137.7 217.3 138.5 216.5 ;
      RECT  135.7 224.3 136.5 223.5 ;
      RECT  139.7 224.3 140.5 223.5 ;
      RECT  136.7 222.8 137.5 222.0 ;
      RECT  138.7 220.0 139.5 219.2 ;
      RECT  141.2 218.6 141.8 218.0 ;
      RECT  134.5 215.5 143.1 214.9 ;
      RECT  134.5 225.9 143.1 225.3 ;
      RECT  146.3 217.3 147.1 216.5 ;
      RECT  144.3 217.3 145.1 216.5 ;
      RECT  146.3 224.7 147.1 223.9 ;
      RECT  144.3 224.7 145.1 223.9 ;
      RECT  144.7 221.0 145.5 220.2 ;
      RECT  146.7 220.9 147.3 220.3 ;
      RECT  143.1 215.5 149.7 214.9 ;
      RECT  143.1 225.9 149.7 225.3 ;
      RECT  136.7 222.8 137.5 222.0 ;
      RECT  138.7 220.0 139.5 219.2 ;
      RECT  146.7 220.9 147.3 220.3 ;
      RECT  134.5 215.5 149.7 214.9 ;
      RECT  134.5 225.9 149.7 225.3 ;
      RECT  137.7 233.9 138.5 234.7 ;
      RECT  135.7 233.9 136.5 234.7 ;
      RECT  139.7 233.9 140.5 234.7 ;
      RECT  137.7 233.9 138.5 234.7 ;
      RECT  135.7 226.9 136.5 227.7 ;
      RECT  139.7 226.9 140.5 227.7 ;
      RECT  136.7 228.4 137.5 229.2 ;
      RECT  138.7 231.2 139.5 232.0 ;
      RECT  141.2 232.6 141.8 233.2 ;
      RECT  134.5 235.7 143.1 236.3 ;
      RECT  134.5 225.3 143.1 225.9 ;
      RECT  146.3 233.9 147.1 234.7 ;
      RECT  144.3 233.9 145.1 234.7 ;
      RECT  146.3 226.5 147.1 227.3 ;
      RECT  144.3 226.5 145.1 227.3 ;
      RECT  144.7 230.2 145.5 231.0 ;
      RECT  146.7 230.3 147.3 230.9 ;
      RECT  143.1 235.7 149.7 236.3 ;
      RECT  143.1 225.3 149.7 225.9 ;
      RECT  136.7 228.4 137.5 229.2 ;
      RECT  138.7 231.2 139.5 232.0 ;
      RECT  146.7 230.3 147.3 230.9 ;
      RECT  134.5 235.7 149.7 236.3 ;
      RECT  134.5 225.3 149.7 225.9 ;
      RECT  137.7 238.1 138.5 237.3 ;
      RECT  135.7 238.1 136.5 237.3 ;
      RECT  139.7 238.1 140.5 237.3 ;
      RECT  137.7 238.1 138.5 237.3 ;
      RECT  135.7 245.1 136.5 244.3 ;
      RECT  139.7 245.1 140.5 244.3 ;
      RECT  136.7 243.6 137.5 242.8 ;
      RECT  138.7 240.8 139.5 240.0 ;
      RECT  141.2 239.4 141.8 238.8 ;
      RECT  134.5 236.3 143.1 235.7 ;
      RECT  134.5 246.7 143.1 246.1 ;
      RECT  146.3 238.1 147.1 237.3 ;
      RECT  144.3 238.1 145.1 237.3 ;
      RECT  146.3 245.5 147.1 244.7 ;
      RECT  144.3 245.5 145.1 244.7 ;
      RECT  144.7 241.8 145.5 241.0 ;
      RECT  146.7 241.7 147.3 241.1 ;
      RECT  143.1 236.3 149.7 235.7 ;
      RECT  143.1 246.7 149.7 246.1 ;
      RECT  136.7 243.6 137.5 242.8 ;
      RECT  138.7 240.8 139.5 240.0 ;
      RECT  146.7 241.7 147.3 241.1 ;
      RECT  134.5 236.3 149.7 235.7 ;
      RECT  134.5 246.7 149.7 246.1 ;
      RECT  137.7 254.7 138.5 255.5 ;
      RECT  135.7 254.7 136.5 255.5 ;
      RECT  139.7 254.7 140.5 255.5 ;
      RECT  137.7 254.7 138.5 255.5 ;
      RECT  135.7 247.7 136.5 248.5 ;
      RECT  139.7 247.7 140.5 248.5 ;
      RECT  136.7 249.2 137.5 250.0 ;
      RECT  138.7 252.0 139.5 252.8 ;
      RECT  141.2 253.4 141.8 254.0 ;
      RECT  134.5 256.5 143.1 257.1 ;
      RECT  134.5 246.1 143.1 246.7 ;
      RECT  146.3 254.7 147.1 255.5 ;
      RECT  144.3 254.7 145.1 255.5 ;
      RECT  146.3 247.3 147.1 248.1 ;
      RECT  144.3 247.3 145.1 248.1 ;
      RECT  144.7 251.0 145.5 251.8 ;
      RECT  146.7 251.1 147.3 251.7 ;
      RECT  143.1 256.5 149.7 257.1 ;
      RECT  143.1 246.1 149.7 246.7 ;
      RECT  136.7 249.2 137.5 250.0 ;
      RECT  138.7 252.0 139.5 252.8 ;
      RECT  146.7 251.1 147.3 251.7 ;
      RECT  134.5 256.5 149.7 257.1 ;
      RECT  134.5 246.1 149.7 246.7 ;
      RECT  137.7 258.9 138.5 258.1 ;
      RECT  135.7 258.9 136.5 258.1 ;
      RECT  139.7 258.9 140.5 258.1 ;
      RECT  137.7 258.9 138.5 258.1 ;
      RECT  135.7 265.9 136.5 265.1 ;
      RECT  139.7 265.9 140.5 265.1 ;
      RECT  136.7 264.4 137.5 263.6 ;
      RECT  138.7 261.6 139.5 260.8 ;
      RECT  141.2 260.2 141.8 259.6 ;
      RECT  134.5 257.1 143.1 256.5 ;
      RECT  134.5 267.5 143.1 266.9 ;
      RECT  146.3 258.9 147.1 258.1 ;
      RECT  144.3 258.9 145.1 258.1 ;
      RECT  146.3 266.3 147.1 265.5 ;
      RECT  144.3 266.3 145.1 265.5 ;
      RECT  144.7 262.6 145.5 261.8 ;
      RECT  146.7 262.5 147.3 261.9 ;
      RECT  143.1 257.1 149.7 256.5 ;
      RECT  143.1 267.5 149.7 266.9 ;
      RECT  136.7 264.4 137.5 263.6 ;
      RECT  138.7 261.6 139.5 260.8 ;
      RECT  146.7 262.5 147.3 261.9 ;
      RECT  134.5 257.1 149.7 256.5 ;
      RECT  134.5 267.5 149.7 266.9 ;
      RECT  137.7 275.5 138.5 276.3 ;
      RECT  135.7 275.5 136.5 276.3 ;
      RECT  139.7 275.5 140.5 276.3 ;
      RECT  137.7 275.5 138.5 276.3 ;
      RECT  135.7 268.5 136.5 269.3 ;
      RECT  139.7 268.5 140.5 269.3 ;
      RECT  136.7 270.0 137.5 270.8 ;
      RECT  138.7 272.8 139.5 273.6 ;
      RECT  141.2 274.2 141.8 274.8 ;
      RECT  134.5 277.3 143.1 277.9 ;
      RECT  134.5 266.9 143.1 267.5 ;
      RECT  146.3 275.5 147.1 276.3 ;
      RECT  144.3 275.5 145.1 276.3 ;
      RECT  146.3 268.1 147.1 268.9 ;
      RECT  144.3 268.1 145.1 268.9 ;
      RECT  144.7 271.8 145.5 272.6 ;
      RECT  146.7 271.9 147.3 272.5 ;
      RECT  143.1 277.3 149.7 277.9 ;
      RECT  143.1 266.9 149.7 267.5 ;
      RECT  136.7 270.0 137.5 270.8 ;
      RECT  138.7 272.8 139.5 273.6 ;
      RECT  146.7 271.9 147.3 272.5 ;
      RECT  134.5 277.3 149.7 277.9 ;
      RECT  134.5 266.9 149.7 267.5 ;
      RECT  137.7 279.7 138.5 278.9 ;
      RECT  135.7 279.7 136.5 278.9 ;
      RECT  139.7 279.7 140.5 278.9 ;
      RECT  137.7 279.7 138.5 278.9 ;
      RECT  135.7 286.7 136.5 285.9 ;
      RECT  139.7 286.7 140.5 285.9 ;
      RECT  136.7 285.2 137.5 284.4 ;
      RECT  138.7 282.4 139.5 281.6 ;
      RECT  141.2 281.0 141.8 280.4 ;
      RECT  134.5 277.9 143.1 277.3 ;
      RECT  134.5 288.3 143.1 287.7 ;
      RECT  146.3 279.7 147.1 278.9 ;
      RECT  144.3 279.7 145.1 278.9 ;
      RECT  146.3 287.1 147.1 286.3 ;
      RECT  144.3 287.1 145.1 286.3 ;
      RECT  144.7 283.4 145.5 282.6 ;
      RECT  146.7 283.3 147.3 282.7 ;
      RECT  143.1 277.9 149.7 277.3 ;
      RECT  143.1 288.3 149.7 287.7 ;
      RECT  136.7 285.2 137.5 284.4 ;
      RECT  138.7 282.4 139.5 281.6 ;
      RECT  146.7 283.3 147.3 282.7 ;
      RECT  134.5 277.9 149.7 277.3 ;
      RECT  134.5 288.3 149.7 287.7 ;
      RECT  137.7 296.3 138.5 297.1 ;
      RECT  135.7 296.3 136.5 297.1 ;
      RECT  139.7 296.3 140.5 297.1 ;
      RECT  137.7 296.3 138.5 297.1 ;
      RECT  135.7 289.3 136.5 290.1 ;
      RECT  139.7 289.3 140.5 290.1 ;
      RECT  136.7 290.8 137.5 291.6 ;
      RECT  138.7 293.6 139.5 294.4 ;
      RECT  141.2 295.0 141.8 295.6 ;
      RECT  134.5 298.1 143.1 298.7 ;
      RECT  134.5 287.7 143.1 288.3 ;
      RECT  146.3 296.3 147.1 297.1 ;
      RECT  144.3 296.3 145.1 297.1 ;
      RECT  146.3 288.9 147.1 289.7 ;
      RECT  144.3 288.9 145.1 289.7 ;
      RECT  144.7 292.6 145.5 293.4 ;
      RECT  146.7 292.7 147.3 293.3 ;
      RECT  143.1 298.1 149.7 298.7 ;
      RECT  143.1 287.7 149.7 288.3 ;
      RECT  136.7 290.8 137.5 291.6 ;
      RECT  138.7 293.6 139.5 294.4 ;
      RECT  146.7 292.7 147.3 293.3 ;
      RECT  134.5 298.1 149.7 298.7 ;
      RECT  134.5 287.7 149.7 288.3 ;
      RECT  137.7 300.5 138.5 299.7 ;
      RECT  135.7 300.5 136.5 299.7 ;
      RECT  139.7 300.5 140.5 299.7 ;
      RECT  137.7 300.5 138.5 299.7 ;
      RECT  135.7 307.5 136.5 306.7 ;
      RECT  139.7 307.5 140.5 306.7 ;
      RECT  136.7 306.0 137.5 305.2 ;
      RECT  138.7 303.2 139.5 302.4 ;
      RECT  141.2 301.8 141.8 301.2 ;
      RECT  134.5 298.7 143.1 298.1 ;
      RECT  134.5 309.1 143.1 308.5 ;
      RECT  146.3 300.5 147.1 299.7 ;
      RECT  144.3 300.5 145.1 299.7 ;
      RECT  146.3 307.9 147.1 307.1 ;
      RECT  144.3 307.9 145.1 307.1 ;
      RECT  144.7 304.2 145.5 303.4 ;
      RECT  146.7 304.1 147.3 303.5 ;
      RECT  143.1 298.7 149.7 298.1 ;
      RECT  143.1 309.1 149.7 308.5 ;
      RECT  136.7 306.0 137.5 305.2 ;
      RECT  138.7 303.2 139.5 302.4 ;
      RECT  146.7 304.1 147.3 303.5 ;
      RECT  134.5 298.7 149.7 298.1 ;
      RECT  134.5 309.1 149.7 308.5 ;
      RECT  137.7 317.1 138.5 317.9 ;
      RECT  135.7 317.1 136.5 317.9 ;
      RECT  139.7 317.1 140.5 317.9 ;
      RECT  137.7 317.1 138.5 317.9 ;
      RECT  135.7 310.1 136.5 310.9 ;
      RECT  139.7 310.1 140.5 310.9 ;
      RECT  136.7 311.6 137.5 312.4 ;
      RECT  138.7 314.4 139.5 315.2 ;
      RECT  141.2 315.8 141.8 316.4 ;
      RECT  134.5 318.9 143.1 319.5 ;
      RECT  134.5 308.5 143.1 309.1 ;
      RECT  146.3 317.1 147.1 317.9 ;
      RECT  144.3 317.1 145.1 317.9 ;
      RECT  146.3 309.7 147.1 310.5 ;
      RECT  144.3 309.7 145.1 310.5 ;
      RECT  144.7 313.4 145.5 314.2 ;
      RECT  146.7 313.5 147.3 314.1 ;
      RECT  143.1 318.9 149.7 319.5 ;
      RECT  143.1 308.5 149.7 309.1 ;
      RECT  136.7 311.6 137.5 312.4 ;
      RECT  138.7 314.4 139.5 315.2 ;
      RECT  146.7 313.5 147.3 314.1 ;
      RECT  134.5 318.9 149.7 319.5 ;
      RECT  134.5 308.5 149.7 309.1 ;
      RECT  137.7 321.3 138.5 320.5 ;
      RECT  135.7 321.3 136.5 320.5 ;
      RECT  139.7 321.3 140.5 320.5 ;
      RECT  137.7 321.3 138.5 320.5 ;
      RECT  135.7 328.3 136.5 327.5 ;
      RECT  139.7 328.3 140.5 327.5 ;
      RECT  136.7 326.8 137.5 326.0 ;
      RECT  138.7 324.0 139.5 323.2 ;
      RECT  141.2 322.6 141.8 322.0 ;
      RECT  134.5 319.5 143.1 318.9 ;
      RECT  134.5 329.9 143.1 329.3 ;
      RECT  146.3 321.3 147.1 320.5 ;
      RECT  144.3 321.3 145.1 320.5 ;
      RECT  146.3 328.7 147.1 327.9 ;
      RECT  144.3 328.7 145.1 327.9 ;
      RECT  144.7 325.0 145.5 324.2 ;
      RECT  146.7 324.9 147.3 324.3 ;
      RECT  143.1 319.5 149.7 318.9 ;
      RECT  143.1 329.9 149.7 329.3 ;
      RECT  136.7 326.8 137.5 326.0 ;
      RECT  138.7 324.0 139.5 323.2 ;
      RECT  146.7 324.9 147.3 324.3 ;
      RECT  134.5 319.5 149.7 318.9 ;
      RECT  134.5 329.9 149.7 329.3 ;
      RECT  137.7 337.9 138.5 338.7 ;
      RECT  135.7 337.9 136.5 338.7 ;
      RECT  139.7 337.9 140.5 338.7 ;
      RECT  137.7 337.9 138.5 338.7 ;
      RECT  135.7 330.9 136.5 331.7 ;
      RECT  139.7 330.9 140.5 331.7 ;
      RECT  136.7 332.4 137.5 333.2 ;
      RECT  138.7 335.2 139.5 336.0 ;
      RECT  141.2 336.6 141.8 337.2 ;
      RECT  134.5 339.7 143.1 340.3 ;
      RECT  134.5 329.3 143.1 329.9 ;
      RECT  146.3 337.9 147.1 338.7 ;
      RECT  144.3 337.9 145.1 338.7 ;
      RECT  146.3 330.5 147.1 331.3 ;
      RECT  144.3 330.5 145.1 331.3 ;
      RECT  144.7 334.2 145.5 335.0 ;
      RECT  146.7 334.3 147.3 334.9 ;
      RECT  143.1 339.7 149.7 340.3 ;
      RECT  143.1 329.3 149.7 329.9 ;
      RECT  136.7 332.4 137.5 333.2 ;
      RECT  138.7 335.2 139.5 336.0 ;
      RECT  146.7 334.3 147.3 334.9 ;
      RECT  134.5 339.7 149.7 340.3 ;
      RECT  134.5 329.3 149.7 329.9 ;
      RECT  137.7 342.1 138.5 341.3 ;
      RECT  135.7 342.1 136.5 341.3 ;
      RECT  139.7 342.1 140.5 341.3 ;
      RECT  137.7 342.1 138.5 341.3 ;
      RECT  135.7 349.1 136.5 348.3 ;
      RECT  139.7 349.1 140.5 348.3 ;
      RECT  136.7 347.6 137.5 346.8 ;
      RECT  138.7 344.8 139.5 344.0 ;
      RECT  141.2 343.4 141.8 342.8 ;
      RECT  134.5 340.3 143.1 339.7 ;
      RECT  134.5 350.7 143.1 350.1 ;
      RECT  146.3 342.1 147.1 341.3 ;
      RECT  144.3 342.1 145.1 341.3 ;
      RECT  146.3 349.5 147.1 348.7 ;
      RECT  144.3 349.5 145.1 348.7 ;
      RECT  144.7 345.8 145.5 345.0 ;
      RECT  146.7 345.7 147.3 345.1 ;
      RECT  143.1 340.3 149.7 339.7 ;
      RECT  143.1 350.7 149.7 350.1 ;
      RECT  136.7 347.6 137.5 346.8 ;
      RECT  138.7 344.8 139.5 344.0 ;
      RECT  146.7 345.7 147.3 345.1 ;
      RECT  134.5 340.3 149.7 339.7 ;
      RECT  134.5 350.7 149.7 350.1 ;
      RECT  146.7 188.7 147.3 189.3 ;
      RECT  146.7 199.5 147.3 200.1 ;
      RECT  146.7 209.5 147.3 210.1 ;
      RECT  146.7 220.3 147.3 220.9 ;
      RECT  146.7 230.3 147.3 230.9 ;
      RECT  146.7 241.1 147.3 241.7 ;
      RECT  146.7 251.1 147.3 251.7 ;
      RECT  146.7 261.9 147.3 262.5 ;
      RECT  146.7 271.9 147.3 272.5 ;
      RECT  146.7 282.7 147.3 283.3 ;
      RECT  146.7 292.7 147.3 293.3 ;
      RECT  146.7 303.5 147.3 304.1 ;
      RECT  146.7 313.5 147.3 314.1 ;
      RECT  146.7 324.3 147.3 324.9 ;
      RECT  146.7 334.3 147.3 334.9 ;
      RECT  146.7 345.1 147.3 345.7 ;
      RECT  153.5 192.3 154.3 193.1 ;
      RECT  151.5 192.3 152.3 193.1 ;
      RECT  155.5 192.3 156.3 193.1 ;
      RECT  153.5 192.3 154.3 193.1 ;
      RECT  151.5 185.3 152.3 186.1 ;
      RECT  155.5 185.3 156.3 186.1 ;
      RECT  152.5 186.8 153.3 187.6 ;
      RECT  154.5 189.6 155.3 190.4 ;
      RECT  157.0 191.0 157.6 191.6 ;
      RECT  150.3 194.1 158.9 194.7 ;
      RECT  150.3 183.7 158.9 184.3 ;
      RECT  162.1 191.5 162.9 192.3 ;
      RECT  160.1 191.5 160.9 192.3 ;
      RECT  162.1 185.3 162.9 186.1 ;
      RECT  160.1 185.3 160.9 186.1 ;
      RECT  160.5 188.4 161.3 189.2 ;
      RECT  162.5 188.5 163.1 189.1 ;
      RECT  158.9 194.1 165.5 194.7 ;
      RECT  158.9 183.7 165.5 184.3 ;
      RECT  152.5 186.8 153.3 187.6 ;
      RECT  154.5 189.6 155.3 190.4 ;
      RECT  162.5 188.5 163.1 189.1 ;
      RECT  150.3 194.1 165.5 194.7 ;
      RECT  150.3 183.7 165.5 184.3 ;
      RECT  153.5 196.5 154.3 195.7 ;
      RECT  151.5 196.5 152.3 195.7 ;
      RECT  155.5 196.5 156.3 195.7 ;
      RECT  153.5 196.5 154.3 195.7 ;
      RECT  151.5 203.5 152.3 202.7 ;
      RECT  155.5 203.5 156.3 202.7 ;
      RECT  152.5 202.0 153.3 201.2 ;
      RECT  154.5 199.2 155.3 198.4 ;
      RECT  157.0 197.8 157.6 197.2 ;
      RECT  150.3 194.7 158.9 194.1 ;
      RECT  150.3 205.1 158.9 204.5 ;
      RECT  162.1 197.3 162.9 196.5 ;
      RECT  160.1 197.3 160.9 196.5 ;
      RECT  162.1 203.5 162.9 202.7 ;
      RECT  160.1 203.5 160.9 202.7 ;
      RECT  160.5 200.4 161.3 199.6 ;
      RECT  162.5 200.3 163.1 199.7 ;
      RECT  158.9 194.7 165.5 194.1 ;
      RECT  158.9 205.1 165.5 204.5 ;
      RECT  152.5 202.0 153.3 201.2 ;
      RECT  154.5 199.2 155.3 198.4 ;
      RECT  162.5 200.3 163.1 199.7 ;
      RECT  150.3 194.7 165.5 194.1 ;
      RECT  150.3 205.1 165.5 204.5 ;
      RECT  153.5 213.1 154.3 213.9 ;
      RECT  151.5 213.1 152.3 213.9 ;
      RECT  155.5 213.1 156.3 213.9 ;
      RECT  153.5 213.1 154.3 213.9 ;
      RECT  151.5 206.1 152.3 206.9 ;
      RECT  155.5 206.1 156.3 206.9 ;
      RECT  152.5 207.6 153.3 208.4 ;
      RECT  154.5 210.4 155.3 211.2 ;
      RECT  157.0 211.8 157.6 212.4 ;
      RECT  150.3 214.9 158.9 215.5 ;
      RECT  150.3 204.5 158.9 205.1 ;
      RECT  162.1 212.3 162.9 213.1 ;
      RECT  160.1 212.3 160.9 213.1 ;
      RECT  162.1 206.1 162.9 206.9 ;
      RECT  160.1 206.1 160.9 206.9 ;
      RECT  160.5 209.2 161.3 210.0 ;
      RECT  162.5 209.3 163.1 209.9 ;
      RECT  158.9 214.9 165.5 215.5 ;
      RECT  158.9 204.5 165.5 205.1 ;
      RECT  152.5 207.6 153.3 208.4 ;
      RECT  154.5 210.4 155.3 211.2 ;
      RECT  162.5 209.3 163.1 209.9 ;
      RECT  150.3 214.9 165.5 215.5 ;
      RECT  150.3 204.5 165.5 205.1 ;
      RECT  153.5 217.3 154.3 216.5 ;
      RECT  151.5 217.3 152.3 216.5 ;
      RECT  155.5 217.3 156.3 216.5 ;
      RECT  153.5 217.3 154.3 216.5 ;
      RECT  151.5 224.3 152.3 223.5 ;
      RECT  155.5 224.3 156.3 223.5 ;
      RECT  152.5 222.8 153.3 222.0 ;
      RECT  154.5 220.0 155.3 219.2 ;
      RECT  157.0 218.6 157.6 218.0 ;
      RECT  150.3 215.5 158.9 214.9 ;
      RECT  150.3 225.9 158.9 225.3 ;
      RECT  162.1 218.1 162.9 217.3 ;
      RECT  160.1 218.1 160.9 217.3 ;
      RECT  162.1 224.3 162.9 223.5 ;
      RECT  160.1 224.3 160.9 223.5 ;
      RECT  160.5 221.2 161.3 220.4 ;
      RECT  162.5 221.1 163.1 220.5 ;
      RECT  158.9 215.5 165.5 214.9 ;
      RECT  158.9 225.9 165.5 225.3 ;
      RECT  152.5 222.8 153.3 222.0 ;
      RECT  154.5 220.0 155.3 219.2 ;
      RECT  162.5 221.1 163.1 220.5 ;
      RECT  150.3 215.5 165.5 214.9 ;
      RECT  150.3 225.9 165.5 225.3 ;
      RECT  153.5 233.9 154.3 234.7 ;
      RECT  151.5 233.9 152.3 234.7 ;
      RECT  155.5 233.9 156.3 234.7 ;
      RECT  153.5 233.9 154.3 234.7 ;
      RECT  151.5 226.9 152.3 227.7 ;
      RECT  155.5 226.9 156.3 227.7 ;
      RECT  152.5 228.4 153.3 229.2 ;
      RECT  154.5 231.2 155.3 232.0 ;
      RECT  157.0 232.6 157.6 233.2 ;
      RECT  150.3 235.7 158.9 236.3 ;
      RECT  150.3 225.3 158.9 225.9 ;
      RECT  162.1 233.1 162.9 233.9 ;
      RECT  160.1 233.1 160.9 233.9 ;
      RECT  162.1 226.9 162.9 227.7 ;
      RECT  160.1 226.9 160.9 227.7 ;
      RECT  160.5 230.0 161.3 230.8 ;
      RECT  162.5 230.1 163.1 230.7 ;
      RECT  158.9 235.7 165.5 236.3 ;
      RECT  158.9 225.3 165.5 225.9 ;
      RECT  152.5 228.4 153.3 229.2 ;
      RECT  154.5 231.2 155.3 232.0 ;
      RECT  162.5 230.1 163.1 230.7 ;
      RECT  150.3 235.7 165.5 236.3 ;
      RECT  150.3 225.3 165.5 225.9 ;
      RECT  153.5 238.1 154.3 237.3 ;
      RECT  151.5 238.1 152.3 237.3 ;
      RECT  155.5 238.1 156.3 237.3 ;
      RECT  153.5 238.1 154.3 237.3 ;
      RECT  151.5 245.1 152.3 244.3 ;
      RECT  155.5 245.1 156.3 244.3 ;
      RECT  152.5 243.6 153.3 242.8 ;
      RECT  154.5 240.8 155.3 240.0 ;
      RECT  157.0 239.4 157.6 238.8 ;
      RECT  150.3 236.3 158.9 235.7 ;
      RECT  150.3 246.7 158.9 246.1 ;
      RECT  162.1 238.9 162.9 238.1 ;
      RECT  160.1 238.9 160.9 238.1 ;
      RECT  162.1 245.1 162.9 244.3 ;
      RECT  160.1 245.1 160.9 244.3 ;
      RECT  160.5 242.0 161.3 241.2 ;
      RECT  162.5 241.9 163.1 241.3 ;
      RECT  158.9 236.3 165.5 235.7 ;
      RECT  158.9 246.7 165.5 246.1 ;
      RECT  152.5 243.6 153.3 242.8 ;
      RECT  154.5 240.8 155.3 240.0 ;
      RECT  162.5 241.9 163.1 241.3 ;
      RECT  150.3 236.3 165.5 235.7 ;
      RECT  150.3 246.7 165.5 246.1 ;
      RECT  153.5 254.7 154.3 255.5 ;
      RECT  151.5 254.7 152.3 255.5 ;
      RECT  155.5 254.7 156.3 255.5 ;
      RECT  153.5 254.7 154.3 255.5 ;
      RECT  151.5 247.7 152.3 248.5 ;
      RECT  155.5 247.7 156.3 248.5 ;
      RECT  152.5 249.2 153.3 250.0 ;
      RECT  154.5 252.0 155.3 252.8 ;
      RECT  157.0 253.4 157.6 254.0 ;
      RECT  150.3 256.5 158.9 257.1 ;
      RECT  150.3 246.1 158.9 246.7 ;
      RECT  162.1 253.9 162.9 254.7 ;
      RECT  160.1 253.9 160.9 254.7 ;
      RECT  162.1 247.7 162.9 248.5 ;
      RECT  160.1 247.7 160.9 248.5 ;
      RECT  160.5 250.8 161.3 251.6 ;
      RECT  162.5 250.9 163.1 251.5 ;
      RECT  158.9 256.5 165.5 257.1 ;
      RECT  158.9 246.1 165.5 246.7 ;
      RECT  152.5 249.2 153.3 250.0 ;
      RECT  154.5 252.0 155.3 252.8 ;
      RECT  162.5 250.9 163.1 251.5 ;
      RECT  150.3 256.5 165.5 257.1 ;
      RECT  150.3 246.1 165.5 246.7 ;
      RECT  153.5 258.9 154.3 258.1 ;
      RECT  151.5 258.9 152.3 258.1 ;
      RECT  155.5 258.9 156.3 258.1 ;
      RECT  153.5 258.9 154.3 258.1 ;
      RECT  151.5 265.9 152.3 265.1 ;
      RECT  155.5 265.9 156.3 265.1 ;
      RECT  152.5 264.4 153.3 263.6 ;
      RECT  154.5 261.6 155.3 260.8 ;
      RECT  157.0 260.2 157.6 259.6 ;
      RECT  150.3 257.1 158.9 256.5 ;
      RECT  150.3 267.5 158.9 266.9 ;
      RECT  162.1 259.7 162.9 258.9 ;
      RECT  160.1 259.7 160.9 258.9 ;
      RECT  162.1 265.9 162.9 265.1 ;
      RECT  160.1 265.9 160.9 265.1 ;
      RECT  160.5 262.8 161.3 262.0 ;
      RECT  162.5 262.7 163.1 262.1 ;
      RECT  158.9 257.1 165.5 256.5 ;
      RECT  158.9 267.5 165.5 266.9 ;
      RECT  152.5 264.4 153.3 263.6 ;
      RECT  154.5 261.6 155.3 260.8 ;
      RECT  162.5 262.7 163.1 262.1 ;
      RECT  150.3 257.1 165.5 256.5 ;
      RECT  150.3 267.5 165.5 266.9 ;
      RECT  153.5 275.5 154.3 276.3 ;
      RECT  151.5 275.5 152.3 276.3 ;
      RECT  155.5 275.5 156.3 276.3 ;
      RECT  153.5 275.5 154.3 276.3 ;
      RECT  151.5 268.5 152.3 269.3 ;
      RECT  155.5 268.5 156.3 269.3 ;
      RECT  152.5 270.0 153.3 270.8 ;
      RECT  154.5 272.8 155.3 273.6 ;
      RECT  157.0 274.2 157.6 274.8 ;
      RECT  150.3 277.3 158.9 277.9 ;
      RECT  150.3 266.9 158.9 267.5 ;
      RECT  162.1 274.7 162.9 275.5 ;
      RECT  160.1 274.7 160.9 275.5 ;
      RECT  162.1 268.5 162.9 269.3 ;
      RECT  160.1 268.5 160.9 269.3 ;
      RECT  160.5 271.6 161.3 272.4 ;
      RECT  162.5 271.7 163.1 272.3 ;
      RECT  158.9 277.3 165.5 277.9 ;
      RECT  158.9 266.9 165.5 267.5 ;
      RECT  152.5 270.0 153.3 270.8 ;
      RECT  154.5 272.8 155.3 273.6 ;
      RECT  162.5 271.7 163.1 272.3 ;
      RECT  150.3 277.3 165.5 277.9 ;
      RECT  150.3 266.9 165.5 267.5 ;
      RECT  153.5 279.7 154.3 278.9 ;
      RECT  151.5 279.7 152.3 278.9 ;
      RECT  155.5 279.7 156.3 278.9 ;
      RECT  153.5 279.7 154.3 278.9 ;
      RECT  151.5 286.7 152.3 285.9 ;
      RECT  155.5 286.7 156.3 285.9 ;
      RECT  152.5 285.2 153.3 284.4 ;
      RECT  154.5 282.4 155.3 281.6 ;
      RECT  157.0 281.0 157.6 280.4 ;
      RECT  150.3 277.9 158.9 277.3 ;
      RECT  150.3 288.3 158.9 287.7 ;
      RECT  162.1 280.5 162.9 279.7 ;
      RECT  160.1 280.5 160.9 279.7 ;
      RECT  162.1 286.7 162.9 285.9 ;
      RECT  160.1 286.7 160.9 285.9 ;
      RECT  160.5 283.6 161.3 282.8 ;
      RECT  162.5 283.5 163.1 282.9 ;
      RECT  158.9 277.9 165.5 277.3 ;
      RECT  158.9 288.3 165.5 287.7 ;
      RECT  152.5 285.2 153.3 284.4 ;
      RECT  154.5 282.4 155.3 281.6 ;
      RECT  162.5 283.5 163.1 282.9 ;
      RECT  150.3 277.9 165.5 277.3 ;
      RECT  150.3 288.3 165.5 287.7 ;
      RECT  153.5 296.3 154.3 297.1 ;
      RECT  151.5 296.3 152.3 297.1 ;
      RECT  155.5 296.3 156.3 297.1 ;
      RECT  153.5 296.3 154.3 297.1 ;
      RECT  151.5 289.3 152.3 290.1 ;
      RECT  155.5 289.3 156.3 290.1 ;
      RECT  152.5 290.8 153.3 291.6 ;
      RECT  154.5 293.6 155.3 294.4 ;
      RECT  157.0 295.0 157.6 295.6 ;
      RECT  150.3 298.1 158.9 298.7 ;
      RECT  150.3 287.7 158.9 288.3 ;
      RECT  162.1 295.5 162.9 296.3 ;
      RECT  160.1 295.5 160.9 296.3 ;
      RECT  162.1 289.3 162.9 290.1 ;
      RECT  160.1 289.3 160.9 290.1 ;
      RECT  160.5 292.4 161.3 293.2 ;
      RECT  162.5 292.5 163.1 293.1 ;
      RECT  158.9 298.1 165.5 298.7 ;
      RECT  158.9 287.7 165.5 288.3 ;
      RECT  152.5 290.8 153.3 291.6 ;
      RECT  154.5 293.6 155.3 294.4 ;
      RECT  162.5 292.5 163.1 293.1 ;
      RECT  150.3 298.1 165.5 298.7 ;
      RECT  150.3 287.7 165.5 288.3 ;
      RECT  153.5 300.5 154.3 299.7 ;
      RECT  151.5 300.5 152.3 299.7 ;
      RECT  155.5 300.5 156.3 299.7 ;
      RECT  153.5 300.5 154.3 299.7 ;
      RECT  151.5 307.5 152.3 306.7 ;
      RECT  155.5 307.5 156.3 306.7 ;
      RECT  152.5 306.0 153.3 305.2 ;
      RECT  154.5 303.2 155.3 302.4 ;
      RECT  157.0 301.8 157.6 301.2 ;
      RECT  150.3 298.7 158.9 298.1 ;
      RECT  150.3 309.1 158.9 308.5 ;
      RECT  162.1 301.3 162.9 300.5 ;
      RECT  160.1 301.3 160.9 300.5 ;
      RECT  162.1 307.5 162.9 306.7 ;
      RECT  160.1 307.5 160.9 306.7 ;
      RECT  160.5 304.4 161.3 303.6 ;
      RECT  162.5 304.3 163.1 303.7 ;
      RECT  158.9 298.7 165.5 298.1 ;
      RECT  158.9 309.1 165.5 308.5 ;
      RECT  152.5 306.0 153.3 305.2 ;
      RECT  154.5 303.2 155.3 302.4 ;
      RECT  162.5 304.3 163.1 303.7 ;
      RECT  150.3 298.7 165.5 298.1 ;
      RECT  150.3 309.1 165.5 308.5 ;
      RECT  153.5 317.1 154.3 317.9 ;
      RECT  151.5 317.1 152.3 317.9 ;
      RECT  155.5 317.1 156.3 317.9 ;
      RECT  153.5 317.1 154.3 317.9 ;
      RECT  151.5 310.1 152.3 310.9 ;
      RECT  155.5 310.1 156.3 310.9 ;
      RECT  152.5 311.6 153.3 312.4 ;
      RECT  154.5 314.4 155.3 315.2 ;
      RECT  157.0 315.8 157.6 316.4 ;
      RECT  150.3 318.9 158.9 319.5 ;
      RECT  150.3 308.5 158.9 309.1 ;
      RECT  162.1 316.3 162.9 317.1 ;
      RECT  160.1 316.3 160.9 317.1 ;
      RECT  162.1 310.1 162.9 310.9 ;
      RECT  160.1 310.1 160.9 310.9 ;
      RECT  160.5 313.2 161.3 314.0 ;
      RECT  162.5 313.3 163.1 313.9 ;
      RECT  158.9 318.9 165.5 319.5 ;
      RECT  158.9 308.5 165.5 309.1 ;
      RECT  152.5 311.6 153.3 312.4 ;
      RECT  154.5 314.4 155.3 315.2 ;
      RECT  162.5 313.3 163.1 313.9 ;
      RECT  150.3 318.9 165.5 319.5 ;
      RECT  150.3 308.5 165.5 309.1 ;
      RECT  153.5 321.3 154.3 320.5 ;
      RECT  151.5 321.3 152.3 320.5 ;
      RECT  155.5 321.3 156.3 320.5 ;
      RECT  153.5 321.3 154.3 320.5 ;
      RECT  151.5 328.3 152.3 327.5 ;
      RECT  155.5 328.3 156.3 327.5 ;
      RECT  152.5 326.8 153.3 326.0 ;
      RECT  154.5 324.0 155.3 323.2 ;
      RECT  157.0 322.6 157.6 322.0 ;
      RECT  150.3 319.5 158.9 318.9 ;
      RECT  150.3 329.9 158.9 329.3 ;
      RECT  162.1 322.1 162.9 321.3 ;
      RECT  160.1 322.1 160.9 321.3 ;
      RECT  162.1 328.3 162.9 327.5 ;
      RECT  160.1 328.3 160.9 327.5 ;
      RECT  160.5 325.2 161.3 324.4 ;
      RECT  162.5 325.1 163.1 324.5 ;
      RECT  158.9 319.5 165.5 318.9 ;
      RECT  158.9 329.9 165.5 329.3 ;
      RECT  152.5 326.8 153.3 326.0 ;
      RECT  154.5 324.0 155.3 323.2 ;
      RECT  162.5 325.1 163.1 324.5 ;
      RECT  150.3 319.5 165.5 318.9 ;
      RECT  150.3 329.9 165.5 329.3 ;
      RECT  153.5 337.9 154.3 338.7 ;
      RECT  151.5 337.9 152.3 338.7 ;
      RECT  155.5 337.9 156.3 338.7 ;
      RECT  153.5 337.9 154.3 338.7 ;
      RECT  151.5 330.9 152.3 331.7 ;
      RECT  155.5 330.9 156.3 331.7 ;
      RECT  152.5 332.4 153.3 333.2 ;
      RECT  154.5 335.2 155.3 336.0 ;
      RECT  157.0 336.6 157.6 337.2 ;
      RECT  150.3 339.7 158.9 340.3 ;
      RECT  150.3 329.3 158.9 329.9 ;
      RECT  162.1 337.1 162.9 337.9 ;
      RECT  160.1 337.1 160.9 337.9 ;
      RECT  162.1 330.9 162.9 331.7 ;
      RECT  160.1 330.9 160.9 331.7 ;
      RECT  160.5 334.0 161.3 334.8 ;
      RECT  162.5 334.1 163.1 334.7 ;
      RECT  158.9 339.7 165.5 340.3 ;
      RECT  158.9 329.3 165.5 329.9 ;
      RECT  152.5 332.4 153.3 333.2 ;
      RECT  154.5 335.2 155.3 336.0 ;
      RECT  162.5 334.1 163.1 334.7 ;
      RECT  150.3 339.7 165.5 340.3 ;
      RECT  150.3 329.3 165.5 329.9 ;
      RECT  153.5 342.1 154.3 341.3 ;
      RECT  151.5 342.1 152.3 341.3 ;
      RECT  155.5 342.1 156.3 341.3 ;
      RECT  153.5 342.1 154.3 341.3 ;
      RECT  151.5 349.1 152.3 348.3 ;
      RECT  155.5 349.1 156.3 348.3 ;
      RECT  152.5 347.6 153.3 346.8 ;
      RECT  154.5 344.8 155.3 344.0 ;
      RECT  157.0 343.4 157.6 342.8 ;
      RECT  150.3 340.3 158.9 339.7 ;
      RECT  150.3 350.7 158.9 350.1 ;
      RECT  162.1 342.9 162.9 342.1 ;
      RECT  160.1 342.9 160.9 342.1 ;
      RECT  162.1 349.1 162.9 348.3 ;
      RECT  160.1 349.1 160.9 348.3 ;
      RECT  160.5 346.0 161.3 345.2 ;
      RECT  162.5 345.9 163.1 345.3 ;
      RECT  158.9 340.3 165.5 339.7 ;
      RECT  158.9 350.7 165.5 350.1 ;
      RECT  152.5 347.6 153.3 346.8 ;
      RECT  154.5 344.8 155.3 344.0 ;
      RECT  162.5 345.9 163.1 345.3 ;
      RECT  150.3 340.3 165.5 339.7 ;
      RECT  150.3 350.7 165.5 350.1 ;
      RECT  152.5 186.8 153.3 187.6 ;
      RECT  152.5 201.2 153.3 202.0 ;
      RECT  152.5 207.6 153.3 208.4 ;
      RECT  152.5 222.0 153.3 222.8 ;
      RECT  152.5 228.4 153.3 229.2 ;
      RECT  152.5 242.8 153.3 243.6 ;
      RECT  152.5 249.2 153.3 250.0 ;
      RECT  152.5 263.6 153.3 264.4 ;
      RECT  152.5 270.0 153.3 270.8 ;
      RECT  152.5 284.4 153.3 285.2 ;
      RECT  152.5 290.8 153.3 291.6 ;
      RECT  152.5 305.2 153.3 306.0 ;
      RECT  152.5 311.6 153.3 312.4 ;
      RECT  152.5 326.0 153.3 326.8 ;
      RECT  152.5 332.4 153.3 333.2 ;
      RECT  152.5 346.8 153.3 347.6 ;
      RECT  162.5 188.5 163.1 189.1 ;
      RECT  162.5 199.7 163.1 200.3 ;
      RECT  162.5 209.3 163.1 209.9 ;
      RECT  162.5 220.5 163.1 221.1 ;
      RECT  162.5 230.1 163.1 230.7 ;
      RECT  162.5 241.3 163.1 241.9 ;
      RECT  162.5 250.9 163.1 251.5 ;
      RECT  162.5 262.1 163.1 262.7 ;
      RECT  162.5 271.7 163.1 272.3 ;
      RECT  162.5 282.9 163.1 283.5 ;
      RECT  162.5 292.5 163.1 293.1 ;
      RECT  162.5 303.7 163.1 304.3 ;
      RECT  162.5 313.3 163.1 313.9 ;
      RECT  162.5 324.5 163.1 325.1 ;
      RECT  162.5 334.1 163.1 334.7 ;
      RECT  162.5 345.3 163.1 345.9 ;
      RECT  162.5 188.5 163.1 189.1 ;
      RECT  162.5 199.7 163.1 200.3 ;
      RECT  162.5 209.3 163.1 209.9 ;
      RECT  162.5 220.5 163.1 221.1 ;
      RECT  162.5 230.1 163.1 230.7 ;
      RECT  162.5 241.3 163.1 241.9 ;
      RECT  162.5 250.9 163.1 251.5 ;
      RECT  162.5 262.1 163.1 262.7 ;
      RECT  162.5 271.7 163.1 272.3 ;
      RECT  162.5 282.9 163.1 283.5 ;
      RECT  162.5 292.5 163.1 293.1 ;
      RECT  162.5 303.7 163.1 304.3 ;
      RECT  162.5 313.3 163.1 313.9 ;
      RECT  162.5 324.5 163.1 325.1 ;
      RECT  162.5 334.1 163.1 334.7 ;
      RECT  162.5 345.3 163.1 345.9 ;
      RECT  1.2 10.2 11.0 10.4 ;
      RECT  15.4 9.6 19.6 10.2 ;
      RECT  18.8 1.2 19.6 5.6 ;
      RECT  7.8 13.6 11.4 14.2 ;
      RECT  18.8 6.2 19.6 9.6 ;
      RECT  7.8 4.4 8.6 4.6 ;
      RECT  10.4 12.0 12.6 12.6 ;
      RECT  1.2 1.2 2.0 6.0 ;
      RECT  11.8 6.6 12.6 6.8 ;
      RECT  7.8 13.4 8.6 13.6 ;
      RECT  11.8 11.8 12.6 12.0 ;
      RECT  4.4 12.0 5.2 12.2 ;
      RECT  12.4 10.6 14.8 11.2 ;
      RECT  5.0 7.4 5.8 7.6 ;
      RECT  18.8 10.2 19.6 18.8 ;
      RECT  15.8 5.4 16.6 5.6 ;
      RECT  14.0 8.2 17.8 8.8 ;
      RECT  6.2 4.6 6.8 6.8 ;
      RECT  8.2 0.6 9.2 3.2 ;
      RECT  17.2 0.6 18.0 5.0 ;
      RECT  9.0 12.0 9.8 12.2 ;
      RECT  17.0 8.8 17.8 9.0 ;
      RECT  10.0 14.8 10.8 18.8 ;
      RECT  4.4 14.0 5.2 14.8 ;
      RECT  14.0 14.0 14.8 14.8 ;
      RECT  6.2 10.4 11.0 10.8 ;
      RECT  1.2 10.0 7.0 10.2 ;
      RECT  3.4 8.6 8.4 9.2 ;
      RECT  10.6 13.4 11.4 13.6 ;
      RECT  4.4 14.8 6.4 15.4 ;
      RECT  2.8 0.6 3.6 5.2 ;
      RECT  7.8 3.8 10.6 4.4 ;
      RECT  20.4 0.6 21.2 2.0 ;
      RECT  1.2 10.4 2.0 18.8 ;
      RECT  2.8 11.0 3.6 19.4 ;
      RECT  14.2 11.2 14.8 12.2 ;
      RECT  14.0 2.6 15.4 3.2 ;
      RECT  8.4 14.8 9.2 19.4 ;
      RECT  11.6 14.8 12.4 19.4 ;
      RECT  14.2 12.2 15.6 13.0 ;
      RECT  12.4 7.4 13.0 10.6 ;
      RECT  2.0 6.6 3.6 6.8 ;
      RECT  4.4 2.6 6.4 3.2 ;
      RECT  5.6 1.2 6.4 2.6 ;
      RECT  14.2 14.8 15.4 18.8 ;
      RECT  6.0 3.8 6.8 4.6 ;
      RECT  10.4 10.8 11.0 12.0 ;
      RECT  7.6 9.2 8.4 9.4 ;
      RECT  14.0 8.0 14.8 8.2 ;
      RECT  10.0 14.2 10.6 14.8 ;
      RECT  4.4 11.4 9.8 12.0 ;
      RECT  10.0 1.2 10.8 3.2 ;
      RECT  0.0 19.4 21.8 20.6 ;
      RECT  5.6 15.4 6.4 18.8 ;
      RECT  17.2 10.8 18.0 19.4 ;
      RECT  1.2 9.8 6.8 10.0 ;
      RECT  3.4 8.4 4.2 8.6 ;
      RECT  11.6 0.6 12.4 3.2 ;
      RECT  14.2 1.2 15.4 2.6 ;
      RECT  0.0 -0.6 21.8 0.6 ;
      RECT  20.4 17.8 21.2 19.4 ;
      RECT  2.0 6.8 13.0 7.4 ;
      RECT  15.8 5.6 19.6 6.2 ;
      RECT  4.4 3.2 5.2 4.0 ;
      RECT  10.0 3.2 10.6 3.8 ;
      RECT  14.0 3.2 14.8 4.0 ;
      RECT  15.4 9.4 16.2 9.6 ;
      RECT  27.4 17.1 28.2 17.9 ;
      RECT  25.4 17.1 26.2 17.9 ;
      RECT  27.4 1.3 28.2 2.1 ;
      RECT  25.4 1.3 26.2 2.1 ;
      RECT  25.8 9.2 26.6 10.0 ;
      RECT  27.8 9.3 28.4 9.9 ;
      RECT  24.2 19.7 30.8 20.3 ;
      RECT  24.2 -0.3 30.8 0.3 ;
      RECT  34.0 15.5 34.8 16.3 ;
      RECT  32.0 15.5 32.8 16.3 ;
      RECT  34.0 2.1 34.8 2.9 ;
      RECT  32.0 2.1 32.8 2.9 ;
      RECT  32.4 8.8 33.2 9.6 ;
      RECT  34.4 8.9 35.0 9.5 ;
      RECT  30.8 19.7 37.4 20.3 ;
      RECT  30.8 -0.3 37.4 0.3 ;
      RECT  0.0 19.4 37.4 20.6 ;
      RECT  0.0 -0.6 37.4 0.6 ;
      RECT  1.2 29.8 11.0 29.6 ;
      RECT  15.4 30.4 19.6 29.8 ;
      RECT  18.8 38.8 19.6 34.4 ;
      RECT  7.8 26.4 11.4 25.8 ;
      RECT  18.8 33.8 19.6 30.4 ;
      RECT  7.8 35.6 8.6 35.4 ;
      RECT  10.4 28.0 12.6 27.4 ;
      RECT  1.2 38.8 2.0 34.0 ;
      RECT  11.8 33.4 12.6 33.2 ;
      RECT  7.8 26.6 8.6 26.4 ;
      RECT  11.8 28.2 12.6 28.0 ;
      RECT  4.4 28.0 5.2 27.8 ;
      RECT  12.4 29.4 14.8 28.8 ;
      RECT  5.0 32.6 5.8 32.4 ;
      RECT  18.8 29.8 19.6 21.2 ;
      RECT  15.8 34.6 16.6 34.4 ;
      RECT  14.0 31.8 17.8 31.2 ;
      RECT  6.2 35.4 6.8 33.2 ;
      RECT  8.2 39.4 9.2 36.8 ;
      RECT  17.2 39.4 18.0 35.0 ;
      RECT  9.0 28.0 9.8 27.8 ;
      RECT  17.0 31.2 17.8 31.0 ;
      RECT  10.0 25.2 10.8 21.2 ;
      RECT  4.4 26.0 5.2 25.2 ;
      RECT  14.0 26.0 14.8 25.2 ;
      RECT  6.2 29.6 11.0 29.2 ;
      RECT  1.2 30.0 7.0 29.8 ;
      RECT  3.4 31.4 8.4 30.8 ;
      RECT  10.6 26.6 11.4 26.4 ;
      RECT  4.4 25.2 6.4 24.6 ;
      RECT  2.8 39.4 3.6 34.8 ;
      RECT  7.8 36.2 10.6 35.6 ;
      RECT  20.4 39.4 21.2 38.0 ;
      RECT  1.2 29.6 2.0 21.2 ;
      RECT  2.8 29.0 3.6 20.6 ;
      RECT  14.2 28.8 14.8 27.8 ;
      RECT  14.0 37.4 15.4 36.8 ;
      RECT  8.4 25.2 9.2 20.6 ;
      RECT  11.6 25.2 12.4 20.6 ;
      RECT  14.2 27.8 15.6 27.0 ;
      RECT  12.4 32.6 13.0 29.4 ;
      RECT  2.0 33.4 3.6 33.2 ;
      RECT  4.4 37.4 6.4 36.8 ;
      RECT  5.6 38.8 6.4 37.4 ;
      RECT  14.2 25.2 15.4 21.2 ;
      RECT  6.0 36.2 6.8 35.4 ;
      RECT  10.4 29.2 11.0 28.0 ;
      RECT  7.6 30.8 8.4 30.6 ;
      RECT  14.0 32.0 14.8 31.8 ;
      RECT  10.0 25.8 10.6 25.2 ;
      RECT  4.4 28.6 9.8 28.0 ;
      RECT  10.0 38.8 10.8 36.8 ;
      RECT  0.0 20.6 21.8 19.4 ;
      RECT  5.6 24.6 6.4 21.2 ;
      RECT  17.2 29.2 18.0 20.6 ;
      RECT  1.2 30.2 6.8 30.0 ;
      RECT  3.4 31.6 4.2 31.4 ;
      RECT  11.6 39.4 12.4 36.8 ;
      RECT  14.2 38.8 15.4 37.4 ;
      RECT  0.0 40.6 21.8 39.4 ;
      RECT  20.4 22.2 21.2 20.6 ;
      RECT  2.0 33.2 13.0 32.6 ;
      RECT  15.8 34.4 19.6 33.8 ;
      RECT  4.4 36.8 5.2 36.0 ;
      RECT  10.0 36.8 10.6 36.2 ;
      RECT  14.0 36.8 14.8 36.0 ;
      RECT  15.4 30.6 16.2 30.4 ;
      RECT  27.4 22.9 28.2 22.1 ;
      RECT  25.4 22.9 26.2 22.1 ;
      RECT  27.4 38.7 28.2 37.9 ;
      RECT  25.4 38.7 26.2 37.9 ;
      RECT  25.8 30.8 26.6 30.0 ;
      RECT  27.8 30.7 28.4 30.1 ;
      RECT  24.2 20.3 30.8 19.7 ;
      RECT  24.2 40.3 30.8 39.7 ;
      RECT  34.0 24.5 34.8 23.7 ;
      RECT  32.0 24.5 32.8 23.7 ;
      RECT  34.0 37.9 34.8 37.1 ;
      RECT  32.0 37.9 32.8 37.1 ;
      RECT  32.4 31.2 33.2 30.4 ;
      RECT  34.4 31.1 35.0 30.5 ;
      RECT  30.8 20.3 37.4 19.7 ;
      RECT  30.8 40.3 37.4 39.7 ;
      RECT  0.0 20.6 37.4 19.4 ;
      RECT  0.0 40.6 37.4 39.4 ;
      RECT  53.2 17.9 54.0 18.7 ;
      RECT  51.2 17.9 52.0 18.7 ;
      RECT  53.2 0.9 54.0 1.7 ;
      RECT  51.2 0.9 52.0 1.7 ;
      RECT  51.6 9.4 52.4 10.2 ;
      RECT  53.6 9.5 54.2 10.1 ;
      RECT  50.0 19.7 56.6 20.3 ;
      RECT  50.0 -0.3 56.6 0.3 ;
      RECT  59.8 17.1 60.6 17.9 ;
      RECT  57.8 17.1 58.6 17.9 ;
      RECT  59.8 1.3 60.6 2.1 ;
      RECT  57.8 1.3 58.6 2.1 ;
      RECT  58.2 9.2 59.0 10.0 ;
      RECT  60.2 9.3 60.8 9.9 ;
      RECT  56.6 19.7 61.8 20.3 ;
      RECT  56.6 -0.3 61.8 0.3 ;
      RECT  65.0 14.7 65.8 15.5 ;
      RECT  63.0 14.7 63.8 15.5 ;
      RECT  65.0 2.5 65.8 3.3 ;
      RECT  63.0 2.5 63.8 3.3 ;
      RECT  63.4 8.6 64.2 9.4 ;
      RECT  65.4 8.7 66.0 9.3 ;
      RECT  61.8 19.7 67.0 20.3 ;
      RECT  61.8 -0.3 67.0 0.3 ;
      RECT  70.1 13.5 74.1 14.1 ;
      RECT  68.2 14.7 69.0 15.5 ;
      RECT  71.6 14.7 72.4 15.5 ;
      RECT  70.1 3.9 74.1 4.5 ;
      RECT  68.2 2.5 69.0 3.3 ;
      RECT  71.6 2.5 72.4 3.3 ;
      RECT  68.6 8.6 69.4 9.4 ;
      RECT  72.1 8.7 72.7 9.3 ;
      RECT  67.0 19.7 75.6 20.3 ;
      RECT  67.0 -0.3 75.6 0.3 ;
      RECT  51.6 9.4 52.4 10.2 ;
      RECT  72.1 8.7 72.7 9.3 ;
      RECT  50.0 19.7 75.6 20.3 ;
      RECT  50.0 -0.3 75.6 0.3 ;
      RECT  53.2 22.1 54.0 21.3 ;
      RECT  51.2 22.1 52.0 21.3 ;
      RECT  53.2 39.1 54.0 38.3 ;
      RECT  51.2 39.1 52.0 38.3 ;
      RECT  51.6 30.6 52.4 29.8 ;
      RECT  53.6 30.5 54.2 29.9 ;
      RECT  50.0 20.3 56.6 19.7 ;
      RECT  50.0 40.3 56.6 39.7 ;
      RECT  59.8 22.1 60.6 21.3 ;
      RECT  57.8 22.1 58.6 21.3 ;
      RECT  61.8 22.1 62.6 21.3 ;
      RECT  59.8 22.1 60.6 21.3 ;
      RECT  57.8 38.7 58.6 37.9 ;
      RECT  61.8 38.7 62.6 37.9 ;
      RECT  58.8 37.2 59.6 36.4 ;
      RECT  60.8 34.4 61.6 33.6 ;
      RECT  63.3 23.4 63.9 22.8 ;
      RECT  56.6 20.3 64.2 19.7 ;
      RECT  56.6 40.3 64.2 39.7 ;
      RECT  67.3 25.7 71.3 25.1 ;
      RECT  68.8 24.5 69.6 23.7 ;
      RECT  65.4 24.5 66.2 23.7 ;
      RECT  67.3 36.5 71.3 35.9 ;
      RECT  68.8 37.9 69.6 37.1 ;
      RECT  65.4 37.9 66.2 37.1 ;
      RECT  65.8 31.2 66.6 30.4 ;
      RECT  69.3 31.1 69.9 30.5 ;
      RECT  64.2 20.3 74.0 19.7 ;
      RECT  64.2 40.3 74.0 39.7 ;
      RECT  65.8 31.2 66.6 30.4 ;
      RECT  69.3 31.1 69.9 30.5 ;
      RECT  64.2 20.3 74.0 19.7 ;
      RECT  64.2 40.3 74.0 39.7 ;
      RECT  58.8 37.2 59.6 36.4 ;
      RECT  60.8 34.4 61.6 33.6 ;
      RECT  69.3 31.1 69.9 30.5 ;
      RECT  56.6 20.3 74.0 19.7 ;
      RECT  56.6 40.3 74.0 39.7 ;
      RECT  53.2 57.9 54.0 58.7 ;
      RECT  51.2 57.9 52.0 58.7 ;
      RECT  55.2 57.9 56.0 58.7 ;
      RECT  53.2 57.9 54.0 58.7 ;
      RECT  51.2 41.3 52.0 42.1 ;
      RECT  55.2 41.3 56.0 42.1 ;
      RECT  52.2 42.8 53.0 43.6 ;
      RECT  54.2 45.6 55.0 46.4 ;
      RECT  56.7 56.6 57.3 57.2 ;
      RECT  50.0 59.7 57.6 60.3 ;
      RECT  50.0 39.7 57.6 40.3 ;
      RECT  60.7 54.3 64.7 54.9 ;
      RECT  62.2 55.5 63.0 56.3 ;
      RECT  58.8 55.5 59.6 56.3 ;
      RECT  60.7 43.5 64.7 44.1 ;
      RECT  62.2 42.1 63.0 42.9 ;
      RECT  58.8 42.1 59.6 42.9 ;
      RECT  59.2 48.8 60.0 49.6 ;
      RECT  62.7 48.9 63.3 49.5 ;
      RECT  57.6 59.7 67.4 60.3 ;
      RECT  57.6 39.7 67.4 40.3 ;
      RECT  59.2 48.8 60.0 49.6 ;
      RECT  62.7 48.9 63.3 49.5 ;
      RECT  57.6 59.7 67.4 60.3 ;
      RECT  57.6 39.7 67.4 40.3 ;
      RECT  52.2 42.8 53.0 43.6 ;
      RECT  54.2 45.6 55.0 46.4 ;
      RECT  62.7 48.9 63.3 49.5 ;
      RECT  50.0 59.7 67.4 60.3 ;
      RECT  50.0 39.7 67.4 40.3 ;
      RECT  53.2 62.1 54.0 61.3 ;
      RECT  51.2 62.1 52.0 61.3 ;
      RECT  53.2 79.1 54.0 78.3 ;
      RECT  51.2 79.1 52.0 78.3 ;
      RECT  51.6 70.6 52.4 69.8 ;
      RECT  53.6 70.5 54.2 69.9 ;
      RECT  50.0 60.3 56.6 59.7 ;
      RECT  50.0 80.3 56.6 79.7 ;
      RECT  59.8 62.1 60.6 61.3 ;
      RECT  57.8 62.1 58.6 61.3 ;
      RECT  59.8 79.1 60.6 78.3 ;
      RECT  57.8 79.1 58.6 78.3 ;
      RECT  58.2 70.6 59.0 69.8 ;
      RECT  60.2 70.5 60.8 69.9 ;
      RECT  56.6 60.3 61.8 59.7 ;
      RECT  56.6 80.3 61.8 79.7 ;
      RECT  65.0 62.9 65.8 62.1 ;
      RECT  63.0 62.9 63.8 62.1 ;
      RECT  65.0 78.7 65.8 77.9 ;
      RECT  63.0 78.7 63.8 77.9 ;
      RECT  63.4 70.8 64.2 70.0 ;
      RECT  65.4 70.7 66.0 70.1 ;
      RECT  61.8 60.3 67.0 59.7 ;
      RECT  61.8 80.3 67.0 79.7 ;
      RECT  70.2 65.3 71.0 64.5 ;
      RECT  68.2 65.3 69.0 64.5 ;
      RECT  70.2 77.5 71.0 76.7 ;
      RECT  68.2 77.5 69.0 76.7 ;
      RECT  68.6 71.4 69.4 70.6 ;
      RECT  70.6 71.3 71.2 70.7 ;
      RECT  67.0 60.3 72.2 59.7 ;
      RECT  67.0 80.3 72.2 79.7 ;
      RECT  51.6 70.6 52.4 69.8 ;
      RECT  70.6 71.3 71.2 70.7 ;
      RECT  50.0 60.3 72.2 59.7 ;
      RECT  50.0 80.3 72.2 79.7 ;
      RECT  53.2 137.9 54.0 138.7 ;
      RECT  51.2 137.9 52.0 138.7 ;
      RECT  53.2 120.9 54.0 121.7 ;
      RECT  51.2 120.9 52.0 121.7 ;
      RECT  51.6 129.4 52.4 130.2 ;
      RECT  53.6 129.5 54.2 130.1 ;
      RECT  50.0 139.7 56.6 140.3 ;
      RECT  50.0 119.7 56.6 120.3 ;
      RECT  53.2 97.9 54.0 98.7 ;
      RECT  51.2 97.9 52.0 98.7 ;
      RECT  55.2 97.9 56.0 98.7 ;
      RECT  53.2 97.9 54.0 98.7 ;
      RECT  57.2 97.9 58.0 98.7 ;
      RECT  55.2 97.9 56.0 98.7 ;
      RECT  51.2 81.3 52.0 82.1 ;
      RECT  57.2 81.3 58.0 82.1 ;
      RECT  51.8 82.8 52.6 83.6 ;
      RECT  54.2 84.2 55.0 85.0 ;
      RECT  56.6 85.6 57.4 86.4 ;
      RECT  58.7 96.7 59.3 97.3 ;
      RECT  50.0 99.7 59.6 100.3 ;
      RECT  50.0 79.7 59.6 80.3 ;
      RECT  62.6 94.7 63.4 95.5 ;
      RECT  60.8 94.7 61.6 95.5 ;
      RECT  64.4 94.7 65.2 95.5 ;
      RECT  62.6 82.5 63.4 83.3 ;
      RECT  60.8 82.5 61.6 83.3 ;
      RECT  64.4 82.5 65.2 83.3 ;
      RECT  61.2 88.6 62.0 89.4 ;
      RECT  63.0 88.7 63.6 89.3 ;
      RECT  59.6 99.7 67.8 100.3 ;
      RECT  59.6 79.7 67.8 80.3 ;
      RECT  61.2 88.6 62.0 89.4 ;
      RECT  63.0 88.7 63.6 89.3 ;
      RECT  59.6 99.7 67.8 100.3 ;
      RECT  59.6 79.7 67.8 80.3 ;
      RECT  51.8 82.8 52.6 83.6 ;
      RECT  54.2 84.2 55.0 85.0 ;
      RECT  56.6 85.6 57.4 86.4 ;
      RECT  63.0 88.7 63.6 89.3 ;
      RECT  50.0 99.7 67.8 100.3 ;
      RECT  50.0 79.7 67.8 80.3 ;
      RECT  53.2 142.1 54.0 141.3 ;
      RECT  51.2 142.1 52.0 141.3 ;
      RECT  55.2 142.1 56.0 141.3 ;
      RECT  53.2 142.1 54.0 141.3 ;
      RECT  57.2 142.1 58.0 141.3 ;
      RECT  55.2 142.1 56.0 141.3 ;
      RECT  51.2 158.7 52.0 157.9 ;
      RECT  57.2 158.7 58.0 157.9 ;
      RECT  51.8 157.2 52.6 156.4 ;
      RECT  54.2 155.8 55.0 155.0 ;
      RECT  56.6 154.4 57.4 153.6 ;
      RECT  58.7 143.3 59.3 142.7 ;
      RECT  50.0 140.3 59.6 139.7 ;
      RECT  50.0 160.3 59.6 159.7 ;
      RECT  62.8 142.9 63.6 142.1 ;
      RECT  60.8 142.9 61.6 142.1 ;
      RECT  62.8 158.7 63.6 157.9 ;
      RECT  60.8 158.7 61.6 157.9 ;
      RECT  61.2 150.8 62.0 150.0 ;
      RECT  63.2 150.7 63.8 150.1 ;
      RECT  59.6 140.3 66.2 139.7 ;
      RECT  59.6 160.3 66.2 159.7 ;
      RECT  61.2 150.8 62.0 150.0 ;
      RECT  63.2 150.7 63.8 150.1 ;
      RECT  59.6 140.3 66.2 139.7 ;
      RECT  59.6 160.3 66.2 159.7 ;
      RECT  51.8 157.2 52.6 156.4 ;
      RECT  54.2 155.8 55.0 155.0 ;
      RECT  56.6 154.4 57.4 153.6 ;
      RECT  63.2 150.7 63.8 150.1 ;
      RECT  50.0 140.3 66.2 139.7 ;
      RECT  50.0 160.3 66.2 159.7 ;
      RECT  29.8 180.3 29.0 181.1 ;
      RECT  31.8 180.3 31.0 181.1 ;
      RECT  29.8 163.7 29.0 164.5 ;
      RECT  31.8 163.7 31.0 164.5 ;
      RECT  31.4 172.0 30.6 172.8 ;
      RECT  29.4 172.1 28.8 172.7 ;
      RECT  33.0 182.1 26.4 182.7 ;
      RECT  33.0 162.5 26.4 163.1 ;
      RECT  23.2 180.3 22.4 181.1 ;
      RECT  25.2 180.3 24.4 181.1 ;
      RECT  23.2 163.7 22.4 164.5 ;
      RECT  25.2 163.7 24.4 164.5 ;
      RECT  24.8 172.0 24.0 172.8 ;
      RECT  22.8 172.1 22.2 172.7 ;
      RECT  26.4 182.1 19.8 182.7 ;
      RECT  26.4 162.5 19.8 163.1 ;
      RECT  16.6 180.3 15.8 181.1 ;
      RECT  18.6 180.3 17.8 181.1 ;
      RECT  16.6 163.7 15.8 164.5 ;
      RECT  18.6 163.7 17.8 164.5 ;
      RECT  18.2 172.0 17.4 172.8 ;
      RECT  16.2 172.1 15.6 172.7 ;
      RECT  19.8 182.1 13.2 182.7 ;
      RECT  19.8 162.5 13.2 163.1 ;
      RECT  10.0 180.3 9.2 181.1 ;
      RECT  12.0 180.3 11.2 181.1 ;
      RECT  10.0 163.7 9.2 164.5 ;
      RECT  12.0 163.7 11.2 164.5 ;
      RECT  11.6 172.0 10.8 172.8 ;
      RECT  9.6 172.1 9.0 172.7 ;
      RECT  13.2 182.1 6.6 182.7 ;
      RECT  13.2 162.5 6.6 163.1 ;
      RECT  3.4 180.3 2.6 181.1 ;
      RECT  5.4 180.3 4.6 181.1 ;
      RECT  3.4 163.7 2.6 164.5 ;
      RECT  5.4 163.7 4.6 164.5 ;
      RECT  5.0 172.0 4.2 172.8 ;
      RECT  3.0 172.1 2.4 172.7 ;
      RECT  6.6 182.1 0.0 182.7 ;
      RECT  6.6 162.5 0.0 163.1 ;
      RECT  29.8 184.5 29.0 183.7 ;
      RECT  31.8 184.5 31.0 183.7 ;
      RECT  29.8 201.1 29.0 200.3 ;
      RECT  31.8 201.1 31.0 200.3 ;
      RECT  31.4 192.8 30.6 192.0 ;
      RECT  29.4 192.7 28.8 192.1 ;
      RECT  33.0 182.7 26.4 182.1 ;
      RECT  33.0 202.3 26.4 201.7 ;
      RECT  23.2 184.5 22.4 183.7 ;
      RECT  25.2 184.5 24.4 183.7 ;
      RECT  23.2 201.1 22.4 200.3 ;
      RECT  25.2 201.1 24.4 200.3 ;
      RECT  24.8 192.8 24.0 192.0 ;
      RECT  22.8 192.7 22.2 192.1 ;
      RECT  26.4 182.7 19.8 182.1 ;
      RECT  26.4 202.3 19.8 201.7 ;
      RECT  16.6 184.5 15.8 183.7 ;
      RECT  18.6 184.5 17.8 183.7 ;
      RECT  16.6 201.1 15.8 200.3 ;
      RECT  18.6 201.1 17.8 200.3 ;
      RECT  18.2 192.8 17.4 192.0 ;
      RECT  16.2 192.7 15.6 192.1 ;
      RECT  19.8 182.7 13.2 182.1 ;
      RECT  19.8 202.3 13.2 201.7 ;
      RECT  10.0 184.5 9.2 183.7 ;
      RECT  12.0 184.5 11.2 183.7 ;
      RECT  10.0 201.1 9.2 200.3 ;
      RECT  12.0 201.1 11.2 200.3 ;
      RECT  11.6 192.8 10.8 192.0 ;
      RECT  9.6 192.7 9.0 192.1 ;
      RECT  13.2 182.7 6.6 182.1 ;
      RECT  13.2 202.3 6.6 201.7 ;
      RECT  3.4 184.5 2.6 183.7 ;
      RECT  5.4 184.5 4.6 183.7 ;
      RECT  3.4 201.1 2.6 200.3 ;
      RECT  5.4 201.1 4.6 200.3 ;
      RECT  5.0 192.8 4.2 192.0 ;
      RECT  3.0 192.7 2.4 192.1 ;
      RECT  6.6 182.7 0.0 182.1 ;
      RECT  6.6 202.3 0.0 201.7 ;
      RECT  29.8 219.5 29.0 220.3 ;
      RECT  31.8 219.5 31.0 220.3 ;
      RECT  29.8 202.9 29.0 203.7 ;
      RECT  31.8 202.9 31.0 203.7 ;
      RECT  31.4 211.2 30.6 212.0 ;
      RECT  29.4 211.3 28.8 211.9 ;
      RECT  33.0 221.3 26.4 221.9 ;
      RECT  33.0 201.7 26.4 202.3 ;
      RECT  23.2 219.5 22.4 220.3 ;
      RECT  25.2 219.5 24.4 220.3 ;
      RECT  23.2 202.9 22.4 203.7 ;
      RECT  25.2 202.9 24.4 203.7 ;
      RECT  24.8 211.2 24.0 212.0 ;
      RECT  22.8 211.3 22.2 211.9 ;
      RECT  26.4 221.3 19.8 221.9 ;
      RECT  26.4 201.7 19.8 202.3 ;
      RECT  16.6 219.5 15.8 220.3 ;
      RECT  18.6 219.5 17.8 220.3 ;
      RECT  16.6 202.9 15.8 203.7 ;
      RECT  18.6 202.9 17.8 203.7 ;
      RECT  18.2 211.2 17.4 212.0 ;
      RECT  16.2 211.3 15.6 211.9 ;
      RECT  19.8 221.3 13.2 221.9 ;
      RECT  19.8 201.7 13.2 202.3 ;
      RECT  10.0 219.5 9.2 220.3 ;
      RECT  12.0 219.5 11.2 220.3 ;
      RECT  10.0 202.9 9.2 203.7 ;
      RECT  12.0 202.9 11.2 203.7 ;
      RECT  11.6 211.2 10.8 212.0 ;
      RECT  9.6 211.3 9.0 211.9 ;
      RECT  13.2 221.3 6.6 221.9 ;
      RECT  13.2 201.7 6.6 202.3 ;
      RECT  3.4 219.5 2.6 220.3 ;
      RECT  5.4 219.5 4.6 220.3 ;
      RECT  3.4 202.9 2.6 203.7 ;
      RECT  5.4 202.9 4.6 203.7 ;
      RECT  5.0 211.2 4.2 212.0 ;
      RECT  3.0 211.3 2.4 211.9 ;
      RECT  6.6 221.3 0.0 221.9 ;
      RECT  6.6 201.7 0.0 202.3 ;
      RECT  29.8 223.7 29.0 222.9 ;
      RECT  31.8 223.7 31.0 222.9 ;
      RECT  29.8 240.3 29.0 239.5 ;
      RECT  31.8 240.3 31.0 239.5 ;
      RECT  31.4 232.0 30.6 231.2 ;
      RECT  29.4 231.9 28.8 231.3 ;
      RECT  33.0 221.9 26.4 221.3 ;
      RECT  33.0 241.5 26.4 240.9 ;
      RECT  23.2 223.7 22.4 222.9 ;
      RECT  25.2 223.7 24.4 222.9 ;
      RECT  23.2 240.3 22.4 239.5 ;
      RECT  25.2 240.3 24.4 239.5 ;
      RECT  24.8 232.0 24.0 231.2 ;
      RECT  22.8 231.9 22.2 231.3 ;
      RECT  26.4 221.9 19.8 221.3 ;
      RECT  26.4 241.5 19.8 240.9 ;
      RECT  16.6 223.7 15.8 222.9 ;
      RECT  18.6 223.7 17.8 222.9 ;
      RECT  16.6 240.3 15.8 239.5 ;
      RECT  18.6 240.3 17.8 239.5 ;
      RECT  18.2 232.0 17.4 231.2 ;
      RECT  16.2 231.9 15.6 231.3 ;
      RECT  19.8 221.9 13.2 221.3 ;
      RECT  19.8 241.5 13.2 240.9 ;
      RECT  10.0 223.7 9.2 222.9 ;
      RECT  12.0 223.7 11.2 222.9 ;
      RECT  10.0 240.3 9.2 239.5 ;
      RECT  12.0 240.3 11.2 239.5 ;
      RECT  11.6 232.0 10.8 231.2 ;
      RECT  9.6 231.9 9.0 231.3 ;
      RECT  13.2 221.9 6.6 221.3 ;
      RECT  13.2 241.5 6.6 240.9 ;
      RECT  3.4 223.7 2.6 222.9 ;
      RECT  5.4 223.7 4.6 222.9 ;
      RECT  3.4 240.3 2.6 239.5 ;
      RECT  5.4 240.3 4.6 239.5 ;
      RECT  5.0 232.0 4.2 231.2 ;
      RECT  3.0 231.9 2.4 231.3 ;
      RECT  6.6 221.9 0.0 221.3 ;
      RECT  6.6 241.5 0.0 240.9 ;
      RECT  29.8 258.7 29.0 259.5 ;
      RECT  31.8 258.7 31.0 259.5 ;
      RECT  29.8 242.1 29.0 242.9 ;
      RECT  31.8 242.1 31.0 242.9 ;
      RECT  31.4 250.4 30.6 251.2 ;
      RECT  29.4 250.5 28.8 251.1 ;
      RECT  33.0 260.5 26.4 261.1 ;
      RECT  33.0 240.9 26.4 241.5 ;
      RECT  23.2 258.7 22.4 259.5 ;
      RECT  25.2 258.7 24.4 259.5 ;
      RECT  23.2 242.1 22.4 242.9 ;
      RECT  25.2 242.1 24.4 242.9 ;
      RECT  24.8 250.4 24.0 251.2 ;
      RECT  22.8 250.5 22.2 251.1 ;
      RECT  26.4 260.5 19.8 261.1 ;
      RECT  26.4 240.9 19.8 241.5 ;
      RECT  16.6 258.7 15.8 259.5 ;
      RECT  18.6 258.7 17.8 259.5 ;
      RECT  16.6 242.1 15.8 242.9 ;
      RECT  18.6 242.1 17.8 242.9 ;
      RECT  18.2 250.4 17.4 251.2 ;
      RECT  16.2 250.5 15.6 251.1 ;
      RECT  19.8 260.5 13.2 261.1 ;
      RECT  19.8 240.9 13.2 241.5 ;
      RECT  10.0 258.7 9.2 259.5 ;
      RECT  12.0 258.7 11.2 259.5 ;
      RECT  10.0 242.1 9.2 242.9 ;
      RECT  12.0 242.1 11.2 242.9 ;
      RECT  11.6 250.4 10.8 251.2 ;
      RECT  9.6 250.5 9.0 251.1 ;
      RECT  13.2 260.5 6.6 261.1 ;
      RECT  13.2 240.9 6.6 241.5 ;
      RECT  3.4 258.7 2.6 259.5 ;
      RECT  5.4 258.7 4.6 259.5 ;
      RECT  3.4 242.1 2.6 242.9 ;
      RECT  5.4 242.1 4.6 242.9 ;
      RECT  5.0 250.4 4.2 251.2 ;
      RECT  3.0 250.5 2.4 251.1 ;
      RECT  6.6 260.5 0.0 261.1 ;
      RECT  6.6 240.9 0.0 241.5 ;
      RECT  29.8 262.9 29.0 262.1 ;
      RECT  31.8 262.9 31.0 262.1 ;
      RECT  29.8 279.5 29.0 278.7 ;
      RECT  31.8 279.5 31.0 278.7 ;
      RECT  31.4 271.2 30.6 270.4 ;
      RECT  29.4 271.1 28.8 270.5 ;
      RECT  33.0 261.1 26.4 260.5 ;
      RECT  33.0 280.7 26.4 280.1 ;
      RECT  23.2 262.9 22.4 262.1 ;
      RECT  25.2 262.9 24.4 262.1 ;
      RECT  23.2 279.5 22.4 278.7 ;
      RECT  25.2 279.5 24.4 278.7 ;
      RECT  24.8 271.2 24.0 270.4 ;
      RECT  22.8 271.1 22.2 270.5 ;
      RECT  26.4 261.1 19.8 260.5 ;
      RECT  26.4 280.7 19.8 280.1 ;
      RECT  16.6 262.9 15.8 262.1 ;
      RECT  18.6 262.9 17.8 262.1 ;
      RECT  16.6 279.5 15.8 278.7 ;
      RECT  18.6 279.5 17.8 278.7 ;
      RECT  18.2 271.2 17.4 270.4 ;
      RECT  16.2 271.1 15.6 270.5 ;
      RECT  19.8 261.1 13.2 260.5 ;
      RECT  19.8 280.7 13.2 280.1 ;
      RECT  10.0 262.9 9.2 262.1 ;
      RECT  12.0 262.9 11.2 262.1 ;
      RECT  10.0 279.5 9.2 278.7 ;
      RECT  12.0 279.5 11.2 278.7 ;
      RECT  11.6 271.2 10.8 270.4 ;
      RECT  9.6 271.1 9.0 270.5 ;
      RECT  13.2 261.1 6.6 260.5 ;
      RECT  13.2 280.7 6.6 280.1 ;
      RECT  3.4 262.9 2.6 262.1 ;
      RECT  5.4 262.9 4.6 262.1 ;
      RECT  3.4 279.5 2.6 278.7 ;
      RECT  5.4 279.5 4.6 278.7 ;
      RECT  5.0 271.2 4.2 270.4 ;
      RECT  3.0 271.1 2.4 270.5 ;
      RECT  6.6 261.1 0.0 260.5 ;
      RECT  6.6 280.7 0.0 280.1 ;
      RECT  29.8 297.9 29.0 298.7 ;
      RECT  31.8 297.9 31.0 298.7 ;
      RECT  29.8 281.3 29.0 282.1 ;
      RECT  31.8 281.3 31.0 282.1 ;
      RECT  31.4 289.6 30.6 290.4 ;
      RECT  29.4 289.7 28.8 290.3 ;
      RECT  33.0 299.7 26.4 300.3 ;
      RECT  33.0 280.1 26.4 280.7 ;
      RECT  23.2 297.9 22.4 298.7 ;
      RECT  25.2 297.9 24.4 298.7 ;
      RECT  23.2 281.3 22.4 282.1 ;
      RECT  25.2 281.3 24.4 282.1 ;
      RECT  24.8 289.6 24.0 290.4 ;
      RECT  22.8 289.7 22.2 290.3 ;
      RECT  26.4 299.7 19.8 300.3 ;
      RECT  26.4 280.1 19.8 280.7 ;
      RECT  16.6 297.9 15.8 298.7 ;
      RECT  18.6 297.9 17.8 298.7 ;
      RECT  16.6 281.3 15.8 282.1 ;
      RECT  18.6 281.3 17.8 282.1 ;
      RECT  18.2 289.6 17.4 290.4 ;
      RECT  16.2 289.7 15.6 290.3 ;
      RECT  19.8 299.7 13.2 300.3 ;
      RECT  19.8 280.1 13.2 280.7 ;
      RECT  10.0 297.9 9.2 298.7 ;
      RECT  12.0 297.9 11.2 298.7 ;
      RECT  10.0 281.3 9.2 282.1 ;
      RECT  12.0 281.3 11.2 282.1 ;
      RECT  11.6 289.6 10.8 290.4 ;
      RECT  9.6 289.7 9.0 290.3 ;
      RECT  13.2 299.7 6.6 300.3 ;
      RECT  13.2 280.1 6.6 280.7 ;
      RECT  3.4 297.9 2.6 298.7 ;
      RECT  5.4 297.9 4.6 298.7 ;
      RECT  3.4 281.3 2.6 282.1 ;
      RECT  5.4 281.3 4.6 282.1 ;
      RECT  5.0 289.6 4.2 290.4 ;
      RECT  3.0 289.7 2.4 290.3 ;
      RECT  6.6 299.7 0.0 300.3 ;
      RECT  6.6 280.1 0.0 280.7 ;
      RECT  29.8 302.1 29.0 301.3 ;
      RECT  31.8 302.1 31.0 301.3 ;
      RECT  29.8 318.7 29.0 317.9 ;
      RECT  31.8 318.7 31.0 317.9 ;
      RECT  31.4 310.4 30.6 309.6 ;
      RECT  29.4 310.3 28.8 309.7 ;
      RECT  33.0 300.3 26.4 299.7 ;
      RECT  33.0 319.9 26.4 319.3 ;
      RECT  23.2 302.1 22.4 301.3 ;
      RECT  25.2 302.1 24.4 301.3 ;
      RECT  23.2 318.7 22.4 317.9 ;
      RECT  25.2 318.7 24.4 317.9 ;
      RECT  24.8 310.4 24.0 309.6 ;
      RECT  22.8 310.3 22.2 309.7 ;
      RECT  26.4 300.3 19.8 299.7 ;
      RECT  26.4 319.9 19.8 319.3 ;
      RECT  16.6 302.1 15.8 301.3 ;
      RECT  18.6 302.1 17.8 301.3 ;
      RECT  16.6 318.7 15.8 317.9 ;
      RECT  18.6 318.7 17.8 317.9 ;
      RECT  18.2 310.4 17.4 309.6 ;
      RECT  16.2 310.3 15.6 309.7 ;
      RECT  19.8 300.3 13.2 299.7 ;
      RECT  19.8 319.9 13.2 319.3 ;
      RECT  10.0 302.1 9.2 301.3 ;
      RECT  12.0 302.1 11.2 301.3 ;
      RECT  10.0 318.7 9.2 317.9 ;
      RECT  12.0 318.7 11.2 317.9 ;
      RECT  11.6 310.4 10.8 309.6 ;
      RECT  9.6 310.3 9.0 309.7 ;
      RECT  13.2 300.3 6.6 299.7 ;
      RECT  13.2 319.9 6.6 319.3 ;
      RECT  3.4 302.1 2.6 301.3 ;
      RECT  5.4 302.1 4.6 301.3 ;
      RECT  3.4 318.7 2.6 317.9 ;
      RECT  5.4 318.7 4.6 317.9 ;
      RECT  5.0 310.4 4.2 309.6 ;
      RECT  3.0 310.3 2.4 309.7 ;
      RECT  6.6 300.3 0.0 299.7 ;
      RECT  6.6 319.9 0.0 319.3 ;
      RECT  29.8 337.1 29.0 337.9 ;
      RECT  31.8 337.1 31.0 337.9 ;
      RECT  29.8 320.5 29.0 321.3 ;
      RECT  31.8 320.5 31.0 321.3 ;
      RECT  31.4 328.8 30.6 329.6 ;
      RECT  29.4 328.9 28.8 329.5 ;
      RECT  33.0 338.9 26.4 339.5 ;
      RECT  33.0 319.3 26.4 319.9 ;
      RECT  23.2 337.1 22.4 337.9 ;
      RECT  25.2 337.1 24.4 337.9 ;
      RECT  23.2 320.5 22.4 321.3 ;
      RECT  25.2 320.5 24.4 321.3 ;
      RECT  24.8 328.8 24.0 329.6 ;
      RECT  22.8 328.9 22.2 329.5 ;
      RECT  26.4 338.9 19.8 339.5 ;
      RECT  26.4 319.3 19.8 319.9 ;
      RECT  16.6 337.1 15.8 337.9 ;
      RECT  18.6 337.1 17.8 337.9 ;
      RECT  16.6 320.5 15.8 321.3 ;
      RECT  18.6 320.5 17.8 321.3 ;
      RECT  18.2 328.8 17.4 329.6 ;
      RECT  16.2 328.9 15.6 329.5 ;
      RECT  19.8 338.9 13.2 339.5 ;
      RECT  19.8 319.3 13.2 319.9 ;
      RECT  10.0 337.1 9.2 337.9 ;
      RECT  12.0 337.1 11.2 337.9 ;
      RECT  10.0 320.5 9.2 321.3 ;
      RECT  12.0 320.5 11.2 321.3 ;
      RECT  11.6 328.8 10.8 329.6 ;
      RECT  9.6 328.9 9.0 329.5 ;
      RECT  13.2 338.9 6.6 339.5 ;
      RECT  13.2 319.3 6.6 319.9 ;
      RECT  3.4 337.1 2.6 337.9 ;
      RECT  5.4 337.1 4.6 337.9 ;
      RECT  3.4 320.5 2.6 321.3 ;
      RECT  5.4 320.5 4.6 321.3 ;
      RECT  5.0 328.8 4.2 329.6 ;
      RECT  3.0 328.9 2.4 329.5 ;
      RECT  6.6 338.9 0.0 339.5 ;
      RECT  6.6 319.3 0.0 319.9 ;
      RECT  53.2 102.1 54.0 101.3 ;
      RECT  51.2 102.1 52.0 101.3 ;
      RECT  55.2 102.1 56.0 101.3 ;
      RECT  53.2 102.1 54.0 101.3 ;
      RECT  51.2 118.7 52.0 117.9 ;
      RECT  55.2 118.7 56.0 117.9 ;
      RECT  52.2 117.2 53.0 116.4 ;
      RECT  54.2 114.4 55.0 113.6 ;
      RECT  56.7 103.4 57.3 102.8 ;
      RECT  50.0 100.3 58.6 99.7 ;
      RECT  50.0 120.3 58.6 119.7 ;
      RECT  61.8 102.1 62.6 101.3 ;
      RECT  59.8 102.1 60.6 101.3 ;
      RECT  61.8 119.1 62.6 118.3 ;
      RECT  59.8 119.1 60.6 118.3 ;
      RECT  60.2 110.6 61.0 109.8 ;
      RECT  62.2 110.5 62.8 109.9 ;
      RECT  58.6 100.3 65.2 99.7 ;
      RECT  58.6 120.3 65.2 119.7 ;
      RECT  68.4 102.1 69.2 101.3 ;
      RECT  66.4 102.1 67.2 101.3 ;
      RECT  68.4 119.1 69.2 118.3 ;
      RECT  66.4 119.1 67.2 118.3 ;
      RECT  66.8 110.6 67.6 109.8 ;
      RECT  68.8 110.5 69.4 109.9 ;
      RECT  65.2 100.3 70.4 99.7 ;
      RECT  65.2 120.3 70.4 119.7 ;
      RECT  60.2 110.6 61.0 109.8 ;
      RECT  68.8 110.5 69.4 109.9 ;
      RECT  58.6 100.3 70.4 99.7 ;
      RECT  58.6 120.3 70.4 119.7 ;
      RECT  56.4 352.2 66.2 352.4 ;
      RECT  70.6 351.6 74.8 352.2 ;
      RECT  74.0 343.2 74.8 347.6 ;
      RECT  63.0 355.6 66.6 356.2 ;
      RECT  74.0 348.2 74.8 351.6 ;
      RECT  63.0 346.4 63.8 346.6 ;
      RECT  65.6 354.0 67.8 354.6 ;
      RECT  56.4 343.2 57.2 348.0 ;
      RECT  67.0 348.6 67.8 348.8 ;
      RECT  63.0 355.4 63.8 355.6 ;
      RECT  67.0 353.8 67.8 354.0 ;
      RECT  59.6 354.0 60.4 354.2 ;
      RECT  67.6 352.6 70.0 353.2 ;
      RECT  60.2 349.4 61.0 349.6 ;
      RECT  74.0 352.2 74.8 360.8 ;
      RECT  71.0 347.4 71.8 347.6 ;
      RECT  69.2 350.2 73.0 350.8 ;
      RECT  61.4 346.6 62.0 348.8 ;
      RECT  63.4 342.6 64.4 345.2 ;
      RECT  72.4 342.6 73.2 347.0 ;
      RECT  64.2 354.0 65.0 354.2 ;
      RECT  72.2 350.8 73.0 351.0 ;
      RECT  65.2 356.8 66.0 360.8 ;
      RECT  59.6 356.0 60.4 356.8 ;
      RECT  69.2 356.0 70.0 356.8 ;
      RECT  61.4 352.4 66.2 352.8 ;
      RECT  56.4 352.0 62.2 352.2 ;
      RECT  58.6 350.6 63.6 351.2 ;
      RECT  65.8 355.4 66.6 355.6 ;
      RECT  59.6 356.8 61.6 357.4 ;
      RECT  58.0 342.6 58.8 347.2 ;
      RECT  63.0 345.8 65.8 346.4 ;
      RECT  75.6 342.6 76.4 344.0 ;
      RECT  56.4 352.4 57.2 360.8 ;
      RECT  58.0 353.0 58.8 361.4 ;
      RECT  69.4 353.2 70.0 354.2 ;
      RECT  69.2 344.6 70.6 345.2 ;
      RECT  63.6 356.8 64.4 361.4 ;
      RECT  66.8 356.8 67.6 361.4 ;
      RECT  69.4 354.2 70.8 355.0 ;
      RECT  67.6 349.4 68.2 352.6 ;
      RECT  57.2 348.6 58.8 348.8 ;
      RECT  59.6 344.6 61.6 345.2 ;
      RECT  60.8 343.2 61.6 344.6 ;
      RECT  69.4 356.8 70.6 360.8 ;
      RECT  61.2 345.8 62.0 346.6 ;
      RECT  65.6 352.8 66.2 354.0 ;
      RECT  62.8 351.2 63.6 351.4 ;
      RECT  69.2 350.0 70.0 350.2 ;
      RECT  65.2 356.2 65.8 356.8 ;
      RECT  59.6 353.4 65.0 354.0 ;
      RECT  65.2 343.2 66.0 345.2 ;
      RECT  55.2 361.4 77.0 362.6 ;
      RECT  60.8 357.4 61.6 360.8 ;
      RECT  72.4 352.8 73.2 361.4 ;
      RECT  56.4 351.8 62.0 352.0 ;
      RECT  58.6 350.4 59.4 350.6 ;
      RECT  66.8 342.6 67.6 345.2 ;
      RECT  69.4 343.2 70.6 344.6 ;
      RECT  55.2 341.4 77.0 342.6 ;
      RECT  75.6 359.8 76.4 361.4 ;
      RECT  57.2 348.8 68.2 349.4 ;
      RECT  71.0 347.6 74.8 348.2 ;
      RECT  59.6 345.2 60.4 346.0 ;
      RECT  65.2 345.2 65.8 345.8 ;
      RECT  69.2 345.2 70.0 346.0 ;
      RECT  70.6 351.4 71.4 351.6 ;
      RECT  56.4 371.8 66.2 371.6 ;
      RECT  70.6 372.4 74.8 371.8 ;
      RECT  74.0 380.8 74.8 376.4 ;
      RECT  63.0 368.4 66.6 367.8 ;
      RECT  74.0 375.8 74.8 372.4 ;
      RECT  63.0 377.6 63.8 377.4 ;
      RECT  65.6 370.0 67.8 369.4 ;
      RECT  56.4 380.8 57.2 376.0 ;
      RECT  67.0 375.4 67.8 375.2 ;
      RECT  63.0 368.6 63.8 368.4 ;
      RECT  67.0 370.2 67.8 370.0 ;
      RECT  59.6 370.0 60.4 369.8 ;
      RECT  67.6 371.4 70.0 370.8 ;
      RECT  60.2 374.6 61.0 374.4 ;
      RECT  74.0 371.8 74.8 363.2 ;
      RECT  71.0 376.6 71.8 376.4 ;
      RECT  69.2 373.8 73.0 373.2 ;
      RECT  61.4 377.4 62.0 375.2 ;
      RECT  63.4 381.4 64.4 378.8 ;
      RECT  72.4 381.4 73.2 377.0 ;
      RECT  64.2 370.0 65.0 369.8 ;
      RECT  72.2 373.2 73.0 373.0 ;
      RECT  65.2 367.2 66.0 363.2 ;
      RECT  59.6 368.0 60.4 367.2 ;
      RECT  69.2 368.0 70.0 367.2 ;
      RECT  61.4 371.6 66.2 371.2 ;
      RECT  56.4 372.0 62.2 371.8 ;
      RECT  58.6 373.4 63.6 372.8 ;
      RECT  65.8 368.6 66.6 368.4 ;
      RECT  59.6 367.2 61.6 366.6 ;
      RECT  58.0 381.4 58.8 376.8 ;
      RECT  63.0 378.2 65.8 377.6 ;
      RECT  75.6 381.4 76.4 380.0 ;
      RECT  56.4 371.6 57.2 363.2 ;
      RECT  58.0 371.0 58.8 362.6 ;
      RECT  69.4 370.8 70.0 369.8 ;
      RECT  69.2 379.4 70.6 378.8 ;
      RECT  63.6 367.2 64.4 362.6 ;
      RECT  66.8 367.2 67.6 362.6 ;
      RECT  69.4 369.8 70.8 369.0 ;
      RECT  67.6 374.6 68.2 371.4 ;
      RECT  57.2 375.4 58.8 375.2 ;
      RECT  59.6 379.4 61.6 378.8 ;
      RECT  60.8 380.8 61.6 379.4 ;
      RECT  69.4 367.2 70.6 363.2 ;
      RECT  61.2 378.2 62.0 377.4 ;
      RECT  65.6 371.2 66.2 370.0 ;
      RECT  62.8 372.8 63.6 372.6 ;
      RECT  69.2 374.0 70.0 373.8 ;
      RECT  65.2 367.8 65.8 367.2 ;
      RECT  59.6 370.6 65.0 370.0 ;
      RECT  65.2 380.8 66.0 378.8 ;
      RECT  55.2 362.6 77.0 361.4 ;
      RECT  60.8 366.6 61.6 363.2 ;
      RECT  72.4 371.2 73.2 362.6 ;
      RECT  56.4 372.2 62.0 372.0 ;
      RECT  58.6 373.6 59.4 373.4 ;
      RECT  66.8 381.4 67.6 378.8 ;
      RECT  69.4 380.8 70.6 379.4 ;
      RECT  55.2 382.6 77.0 381.4 ;
      RECT  75.6 364.2 76.4 362.6 ;
      RECT  57.2 375.2 68.2 374.6 ;
      RECT  71.0 376.4 74.8 375.8 ;
      RECT  59.6 378.8 60.4 378.0 ;
      RECT  65.2 378.8 65.8 378.2 ;
      RECT  69.2 378.8 70.0 378.0 ;
      RECT  70.6 372.6 71.4 372.4 ;
      RECT  56.4 392.2 66.2 392.4 ;
      RECT  70.6 391.6 74.8 392.2 ;
      RECT  74.0 383.2 74.8 387.6 ;
      RECT  63.0 395.6 66.6 396.2 ;
      RECT  74.0 388.2 74.8 391.6 ;
      RECT  63.0 386.4 63.8 386.6 ;
      RECT  65.6 394.0 67.8 394.6 ;
      RECT  56.4 383.2 57.2 388.0 ;
      RECT  67.0 388.6 67.8 388.8 ;
      RECT  63.0 395.4 63.8 395.6 ;
      RECT  67.0 393.8 67.8 394.0 ;
      RECT  59.6 394.0 60.4 394.2 ;
      RECT  67.6 392.6 70.0 393.2 ;
      RECT  60.2 389.4 61.0 389.6 ;
      RECT  74.0 392.2 74.8 400.8 ;
      RECT  71.0 387.4 71.8 387.6 ;
      RECT  69.2 390.2 73.0 390.8 ;
      RECT  61.4 386.6 62.0 388.8 ;
      RECT  63.4 382.6 64.4 385.2 ;
      RECT  72.4 382.6 73.2 387.0 ;
      RECT  64.2 394.0 65.0 394.2 ;
      RECT  72.2 390.8 73.0 391.0 ;
      RECT  65.2 396.8 66.0 400.8 ;
      RECT  59.6 396.0 60.4 396.8 ;
      RECT  69.2 396.0 70.0 396.8 ;
      RECT  61.4 392.4 66.2 392.8 ;
      RECT  56.4 392.0 62.2 392.2 ;
      RECT  58.6 390.6 63.6 391.2 ;
      RECT  65.8 395.4 66.6 395.6 ;
      RECT  59.6 396.8 61.6 397.4 ;
      RECT  58.0 382.6 58.8 387.2 ;
      RECT  63.0 385.8 65.8 386.4 ;
      RECT  75.6 382.6 76.4 384.0 ;
      RECT  56.4 392.4 57.2 400.8 ;
      RECT  58.0 393.0 58.8 401.4 ;
      RECT  69.4 393.2 70.0 394.2 ;
      RECT  69.2 384.6 70.6 385.2 ;
      RECT  63.6 396.8 64.4 401.4 ;
      RECT  66.8 396.8 67.6 401.4 ;
      RECT  69.4 394.2 70.8 395.0 ;
      RECT  67.6 389.4 68.2 392.6 ;
      RECT  57.2 388.6 58.8 388.8 ;
      RECT  59.6 384.6 61.6 385.2 ;
      RECT  60.8 383.2 61.6 384.6 ;
      RECT  69.4 396.8 70.6 400.8 ;
      RECT  61.2 385.8 62.0 386.6 ;
      RECT  65.6 392.8 66.2 394.0 ;
      RECT  62.8 391.2 63.6 391.4 ;
      RECT  69.2 390.0 70.0 390.2 ;
      RECT  65.2 396.2 65.8 396.8 ;
      RECT  59.6 393.4 65.0 394.0 ;
      RECT  65.2 383.2 66.0 385.2 ;
      RECT  55.2 401.4 77.0 402.6 ;
      RECT  60.8 397.4 61.6 400.8 ;
      RECT  72.4 392.8 73.2 401.4 ;
      RECT  56.4 391.8 62.0 392.0 ;
      RECT  58.6 390.4 59.4 390.6 ;
      RECT  66.8 382.6 67.6 385.2 ;
      RECT  69.4 383.2 70.6 384.6 ;
      RECT  55.2 381.4 77.0 382.6 ;
      RECT  75.6 399.8 76.4 401.4 ;
      RECT  57.2 388.8 68.2 389.4 ;
      RECT  71.0 387.6 74.8 388.2 ;
      RECT  59.6 385.2 60.4 386.0 ;
      RECT  65.2 385.2 65.8 385.8 ;
      RECT  69.2 385.2 70.0 386.0 ;
      RECT  70.6 391.4 71.4 391.6 ;
      RECT  56.4 411.8 66.2 411.6 ;
      RECT  70.6 412.4 74.8 411.8 ;
      RECT  74.0 420.8 74.8 416.4 ;
      RECT  63.0 408.4 66.6 407.8 ;
      RECT  74.0 415.8 74.8 412.4 ;
      RECT  63.0 417.6 63.8 417.4 ;
      RECT  65.6 410.0 67.8 409.4 ;
      RECT  56.4 420.8 57.2 416.0 ;
      RECT  67.0 415.4 67.8 415.2 ;
      RECT  63.0 408.6 63.8 408.4 ;
      RECT  67.0 410.2 67.8 410.0 ;
      RECT  59.6 410.0 60.4 409.8 ;
      RECT  67.6 411.4 70.0 410.8 ;
      RECT  60.2 414.6 61.0 414.4 ;
      RECT  74.0 411.8 74.8 403.2 ;
      RECT  71.0 416.6 71.8 416.4 ;
      RECT  69.2 413.8 73.0 413.2 ;
      RECT  61.4 417.4 62.0 415.2 ;
      RECT  63.4 421.4 64.4 418.8 ;
      RECT  72.4 421.4 73.2 417.0 ;
      RECT  64.2 410.0 65.0 409.8 ;
      RECT  72.2 413.2 73.0 413.0 ;
      RECT  65.2 407.2 66.0 403.2 ;
      RECT  59.6 408.0 60.4 407.2 ;
      RECT  69.2 408.0 70.0 407.2 ;
      RECT  61.4 411.6 66.2 411.2 ;
      RECT  56.4 412.0 62.2 411.8 ;
      RECT  58.6 413.4 63.6 412.8 ;
      RECT  65.8 408.6 66.6 408.4 ;
      RECT  59.6 407.2 61.6 406.6 ;
      RECT  58.0 421.4 58.8 416.8 ;
      RECT  63.0 418.2 65.8 417.6 ;
      RECT  75.6 421.4 76.4 420.0 ;
      RECT  56.4 411.6 57.2 403.2 ;
      RECT  58.0 411.0 58.8 402.6 ;
      RECT  69.4 410.8 70.0 409.8 ;
      RECT  69.2 419.4 70.6 418.8 ;
      RECT  63.6 407.2 64.4 402.6 ;
      RECT  66.8 407.2 67.6 402.6 ;
      RECT  69.4 409.8 70.8 409.0 ;
      RECT  67.6 414.6 68.2 411.4 ;
      RECT  57.2 415.4 58.8 415.2 ;
      RECT  59.6 419.4 61.6 418.8 ;
      RECT  60.8 420.8 61.6 419.4 ;
      RECT  69.4 407.2 70.6 403.2 ;
      RECT  61.2 418.2 62.0 417.4 ;
      RECT  65.6 411.2 66.2 410.0 ;
      RECT  62.8 412.8 63.6 412.6 ;
      RECT  69.2 414.0 70.0 413.8 ;
      RECT  65.2 407.8 65.8 407.2 ;
      RECT  59.6 410.6 65.0 410.0 ;
      RECT  65.2 420.8 66.0 418.8 ;
      RECT  55.2 402.6 77.0 401.4 ;
      RECT  60.8 406.6 61.6 403.2 ;
      RECT  72.4 411.2 73.2 402.6 ;
      RECT  56.4 412.2 62.0 412.0 ;
      RECT  58.6 413.6 59.4 413.4 ;
      RECT  66.8 421.4 67.6 418.8 ;
      RECT  69.4 420.8 70.6 419.4 ;
      RECT  55.2 422.6 77.0 421.4 ;
      RECT  75.6 404.2 76.4 402.6 ;
      RECT  57.2 415.2 68.2 414.6 ;
      RECT  71.0 416.4 74.8 415.8 ;
      RECT  59.6 418.8 60.4 418.0 ;
      RECT  65.2 418.8 65.8 418.2 ;
      RECT  69.2 418.8 70.0 418.0 ;
      RECT  70.6 412.6 71.4 412.4 ;
      RECT  100.0 41.2 109.8 41.4 ;
      RECT  114.2 40.6 118.4 41.2 ;
      RECT  117.6 32.2 118.4 36.6 ;
      RECT  106.6 44.6 110.2 45.2 ;
      RECT  117.6 37.2 118.4 40.6 ;
      RECT  106.6 35.4 107.4 35.6 ;
      RECT  109.2 43.0 111.4 43.6 ;
      RECT  100.0 32.2 100.8 37.0 ;
      RECT  110.6 37.6 111.4 37.8 ;
      RECT  106.6 44.4 107.4 44.6 ;
      RECT  110.6 42.8 111.4 43.0 ;
      RECT  103.2 43.0 104.0 43.2 ;
      RECT  111.2 41.6 113.6 42.2 ;
      RECT  103.8 38.4 104.6 38.6 ;
      RECT  117.6 41.2 118.4 49.8 ;
      RECT  114.6 36.4 115.4 36.6 ;
      RECT  112.8 39.2 116.6 39.8 ;
      RECT  105.0 35.6 105.6 37.8 ;
      RECT  107.0 31.6 108.0 34.2 ;
      RECT  116.0 31.6 116.8 36.0 ;
      RECT  107.8 43.0 108.6 43.2 ;
      RECT  115.8 39.8 116.6 40.0 ;
      RECT  108.8 45.8 109.6 49.8 ;
      RECT  103.2 45.0 104.0 45.8 ;
      RECT  112.8 45.0 113.6 45.8 ;
      RECT  105.0 41.4 109.8 41.8 ;
      RECT  100.0 41.0 105.8 41.2 ;
      RECT  102.2 39.6 107.2 40.2 ;
      RECT  109.4 44.4 110.2 44.6 ;
      RECT  103.2 45.8 105.2 46.4 ;
      RECT  101.6 31.6 102.4 36.2 ;
      RECT  106.6 34.8 109.4 35.4 ;
      RECT  119.2 31.6 120.0 33.0 ;
      RECT  100.0 41.4 100.8 49.8 ;
      RECT  101.6 42.0 102.4 50.4 ;
      RECT  113.0 42.2 113.6 43.2 ;
      RECT  112.8 33.6 114.2 34.2 ;
      RECT  107.2 45.8 108.0 50.4 ;
      RECT  110.4 45.8 111.2 50.4 ;
      RECT  113.0 43.2 114.4 44.0 ;
      RECT  111.2 38.4 111.8 41.6 ;
      RECT  100.8 37.6 102.4 37.8 ;
      RECT  103.2 33.6 105.2 34.2 ;
      RECT  104.4 32.2 105.2 33.6 ;
      RECT  113.0 45.8 114.2 49.8 ;
      RECT  104.8 34.8 105.6 35.6 ;
      RECT  109.2 41.8 109.8 43.0 ;
      RECT  106.4 40.2 107.2 40.4 ;
      RECT  112.8 39.0 113.6 39.2 ;
      RECT  108.8 45.2 109.4 45.8 ;
      RECT  103.2 42.4 108.6 43.0 ;
      RECT  108.8 32.2 109.6 34.2 ;
      RECT  98.8 50.4 120.6 51.6 ;
      RECT  104.4 46.4 105.2 49.8 ;
      RECT  116.0 41.8 116.8 50.4 ;
      RECT  100.0 40.8 105.6 41.0 ;
      RECT  102.2 39.4 103.0 39.6 ;
      RECT  110.4 31.6 111.2 34.2 ;
      RECT  113.0 32.2 114.2 33.6 ;
      RECT  98.8 30.4 120.6 31.6 ;
      RECT  119.2 48.8 120.0 50.4 ;
      RECT  100.8 37.8 111.8 38.4 ;
      RECT  114.6 36.6 118.4 37.2 ;
      RECT  103.2 34.2 104.0 35.0 ;
      RECT  108.8 34.2 109.4 34.8 ;
      RECT  112.8 34.2 113.6 35.0 ;
      RECT  114.2 40.4 115.0 40.6 ;
      RECT  121.8 41.2 131.6 41.4 ;
      RECT  136.0 40.6 140.2 41.2 ;
      RECT  139.4 32.2 140.2 36.6 ;
      RECT  128.4 44.6 132.0 45.2 ;
      RECT  139.4 37.2 140.2 40.6 ;
      RECT  128.4 35.4 129.2 35.6 ;
      RECT  131.0 43.0 133.2 43.6 ;
      RECT  121.8 32.2 122.6 37.0 ;
      RECT  132.4 37.6 133.2 37.8 ;
      RECT  128.4 44.4 129.2 44.6 ;
      RECT  132.4 42.8 133.2 43.0 ;
      RECT  125.0 43.0 125.8 43.2 ;
      RECT  133.0 41.6 135.4 42.2 ;
      RECT  125.6 38.4 126.4 38.6 ;
      RECT  139.4 41.2 140.2 49.8 ;
      RECT  136.4 36.4 137.2 36.6 ;
      RECT  134.6 39.2 138.4 39.8 ;
      RECT  126.8 35.6 127.4 37.8 ;
      RECT  128.8 31.6 129.8 34.2 ;
      RECT  137.8 31.6 138.6 36.0 ;
      RECT  129.6 43.0 130.4 43.2 ;
      RECT  137.6 39.8 138.4 40.0 ;
      RECT  130.6 45.8 131.4 49.8 ;
      RECT  125.0 45.0 125.8 45.8 ;
      RECT  134.6 45.0 135.4 45.8 ;
      RECT  126.8 41.4 131.6 41.8 ;
      RECT  121.8 41.0 127.6 41.2 ;
      RECT  124.0 39.6 129.0 40.2 ;
      RECT  131.2 44.4 132.0 44.6 ;
      RECT  125.0 45.8 127.0 46.4 ;
      RECT  123.4 31.6 124.2 36.2 ;
      RECT  128.4 34.8 131.2 35.4 ;
      RECT  141.0 31.6 141.8 33.0 ;
      RECT  121.8 41.4 122.6 49.8 ;
      RECT  123.4 42.0 124.2 50.4 ;
      RECT  134.8 42.2 135.4 43.2 ;
      RECT  134.6 33.6 136.0 34.2 ;
      RECT  129.0 45.8 129.8 50.4 ;
      RECT  132.2 45.8 133.0 50.4 ;
      RECT  134.8 43.2 136.2 44.0 ;
      RECT  133.0 38.4 133.6 41.6 ;
      RECT  122.6 37.6 124.2 37.8 ;
      RECT  125.0 33.6 127.0 34.2 ;
      RECT  126.2 32.2 127.0 33.6 ;
      RECT  134.8 45.8 136.0 49.8 ;
      RECT  126.6 34.8 127.4 35.6 ;
      RECT  131.0 41.8 131.6 43.0 ;
      RECT  128.2 40.2 129.0 40.4 ;
      RECT  134.6 39.0 135.4 39.2 ;
      RECT  130.6 45.2 131.2 45.8 ;
      RECT  125.0 42.4 130.4 43.0 ;
      RECT  130.6 32.2 131.4 34.2 ;
      RECT  120.6 50.4 142.4 51.6 ;
      RECT  126.2 46.4 127.0 49.8 ;
      RECT  137.8 41.8 138.6 50.4 ;
      RECT  121.8 40.8 127.4 41.0 ;
      RECT  124.0 39.4 124.8 39.6 ;
      RECT  132.2 31.6 133.0 34.2 ;
      RECT  134.8 32.2 136.0 33.6 ;
      RECT  120.6 30.4 142.4 31.6 ;
      RECT  141.0 48.8 141.8 50.4 ;
      RECT  122.6 37.8 133.6 38.4 ;
      RECT  136.4 36.6 140.2 37.2 ;
      RECT  125.0 34.2 125.8 35.0 ;
      RECT  130.6 34.2 131.2 34.8 ;
      RECT  134.6 34.2 135.4 35.0 ;
      RECT  136.0 40.4 136.8 40.6 ;
   LAYER  m2 ;
      RECT  184.1 183.6 184.9 194.4 ;
      RECT  187.5 193.6 188.3 194.4 ;
      RECT  189.3 185.2 190.1 194.4 ;
      RECT  185.7 183.6 186.5 194.4 ;
      RECT  190.9 183.6 191.7 194.4 ;
      RECT  188.5 184.4 190.1 185.2 ;
      RECT  189.3 183.6 190.1 184.4 ;
      RECT  184.1 204.4 184.9 193.6 ;
      RECT  187.5 194.4 188.3 193.6 ;
      RECT  189.3 202.8 190.1 193.6 ;
      RECT  185.7 204.4 186.5 193.6 ;
      RECT  190.9 204.4 191.7 193.6 ;
      RECT  188.5 203.6 190.1 202.8 ;
      RECT  189.3 204.4 190.1 203.6 ;
      RECT  184.1 204.4 184.9 215.2 ;
      RECT  187.5 214.4 188.3 215.2 ;
      RECT  189.3 206.0 190.1 215.2 ;
      RECT  185.7 204.4 186.5 215.2 ;
      RECT  190.9 204.4 191.7 215.2 ;
      RECT  188.5 205.2 190.1 206.0 ;
      RECT  189.3 204.4 190.1 205.2 ;
      RECT  184.1 225.2 184.9 214.4 ;
      RECT  187.5 215.2 188.3 214.4 ;
      RECT  189.3 223.6 190.1 214.4 ;
      RECT  185.7 225.2 186.5 214.4 ;
      RECT  190.9 225.2 191.7 214.4 ;
      RECT  188.5 224.4 190.1 223.6 ;
      RECT  189.3 225.2 190.1 224.4 ;
      RECT  184.1 225.2 184.9 236.0 ;
      RECT  187.5 235.2 188.3 236.0 ;
      RECT  189.3 226.8 190.1 236.0 ;
      RECT  185.7 225.2 186.5 236.0 ;
      RECT  190.9 225.2 191.7 236.0 ;
      RECT  188.5 226.0 190.1 226.8 ;
      RECT  189.3 225.2 190.1 226.0 ;
      RECT  184.1 246.0 184.9 235.2 ;
      RECT  187.5 236.0 188.3 235.2 ;
      RECT  189.3 244.4 190.1 235.2 ;
      RECT  185.7 246.0 186.5 235.2 ;
      RECT  190.9 246.0 191.7 235.2 ;
      RECT  188.5 245.2 190.1 244.4 ;
      RECT  189.3 246.0 190.1 245.2 ;
      RECT  184.1 246.0 184.9 256.8 ;
      RECT  187.5 256.0 188.3 256.8 ;
      RECT  189.3 247.6 190.1 256.8 ;
      RECT  185.7 246.0 186.5 256.8 ;
      RECT  190.9 246.0 191.7 256.8 ;
      RECT  188.5 246.8 190.1 247.6 ;
      RECT  189.3 246.0 190.1 246.8 ;
      RECT  184.1 266.8 184.9 256.0 ;
      RECT  187.5 256.8 188.3 256.0 ;
      RECT  189.3 265.2 190.1 256.0 ;
      RECT  185.7 266.8 186.5 256.0 ;
      RECT  190.9 266.8 191.7 256.0 ;
      RECT  188.5 266.0 190.1 265.2 ;
      RECT  189.3 266.8 190.1 266.0 ;
      RECT  184.1 266.8 184.9 277.6 ;
      RECT  187.5 276.8 188.3 277.6 ;
      RECT  189.3 268.4 190.1 277.6 ;
      RECT  185.7 266.8 186.5 277.6 ;
      RECT  190.9 266.8 191.7 277.6 ;
      RECT  188.5 267.6 190.1 268.4 ;
      RECT  189.3 266.8 190.1 267.6 ;
      RECT  184.1 287.6 184.9 276.8 ;
      RECT  187.5 277.6 188.3 276.8 ;
      RECT  189.3 286.0 190.1 276.8 ;
      RECT  185.7 287.6 186.5 276.8 ;
      RECT  190.9 287.6 191.7 276.8 ;
      RECT  188.5 286.8 190.1 286.0 ;
      RECT  189.3 287.6 190.1 286.8 ;
      RECT  184.1 287.6 184.9 298.4 ;
      RECT  187.5 297.6 188.3 298.4 ;
      RECT  189.3 289.2 190.1 298.4 ;
      RECT  185.7 287.6 186.5 298.4 ;
      RECT  190.9 287.6 191.7 298.4 ;
      RECT  188.5 288.4 190.1 289.2 ;
      RECT  189.3 287.6 190.1 288.4 ;
      RECT  184.1 308.4 184.9 297.6 ;
      RECT  187.5 298.4 188.3 297.6 ;
      RECT  189.3 306.8 190.1 297.6 ;
      RECT  185.7 308.4 186.5 297.6 ;
      RECT  190.9 308.4 191.7 297.6 ;
      RECT  188.5 307.6 190.1 306.8 ;
      RECT  189.3 308.4 190.1 307.6 ;
      RECT  184.1 308.4 184.9 319.2 ;
      RECT  187.5 318.4 188.3 319.2 ;
      RECT  189.3 310.0 190.1 319.2 ;
      RECT  185.7 308.4 186.5 319.2 ;
      RECT  190.9 308.4 191.7 319.2 ;
      RECT  188.5 309.2 190.1 310.0 ;
      RECT  189.3 308.4 190.1 309.2 ;
      RECT  184.1 329.2 184.9 318.4 ;
      RECT  187.5 319.2 188.3 318.4 ;
      RECT  189.3 327.6 190.1 318.4 ;
      RECT  185.7 329.2 186.5 318.4 ;
      RECT  190.9 329.2 191.7 318.4 ;
      RECT  188.5 328.4 190.1 327.6 ;
      RECT  189.3 329.2 190.1 328.4 ;
      RECT  184.1 329.2 184.9 340.0 ;
      RECT  187.5 339.2 188.3 340.0 ;
      RECT  189.3 330.8 190.1 340.0 ;
      RECT  185.7 329.2 186.5 340.0 ;
      RECT  190.9 329.2 191.7 340.0 ;
      RECT  188.5 330.0 190.1 330.8 ;
      RECT  189.3 329.2 190.1 330.0 ;
      RECT  184.1 350.0 184.9 339.2 ;
      RECT  187.5 340.0 188.3 339.2 ;
      RECT  189.3 348.4 190.1 339.2 ;
      RECT  185.7 350.0 186.5 339.2 ;
      RECT  190.9 350.0 191.7 339.2 ;
      RECT  188.5 349.2 190.1 348.4 ;
      RECT  189.3 350.0 190.1 349.2 ;
      RECT  190.9 183.6 191.7 194.4 ;
      RECT  194.3 193.6 195.1 194.4 ;
      RECT  196.1 185.2 196.9 194.4 ;
      RECT  192.5 183.6 193.3 194.4 ;
      RECT  197.7 183.6 198.5 194.4 ;
      RECT  195.3 184.4 196.9 185.2 ;
      RECT  196.1 183.6 196.9 184.4 ;
      RECT  190.9 204.4 191.7 193.6 ;
      RECT  194.3 194.4 195.1 193.6 ;
      RECT  196.1 202.8 196.9 193.6 ;
      RECT  192.5 204.4 193.3 193.6 ;
      RECT  197.7 204.4 198.5 193.6 ;
      RECT  195.3 203.6 196.9 202.8 ;
      RECT  196.1 204.4 196.9 203.6 ;
      RECT  190.9 204.4 191.7 215.2 ;
      RECT  194.3 214.4 195.1 215.2 ;
      RECT  196.1 206.0 196.9 215.2 ;
      RECT  192.5 204.4 193.3 215.2 ;
      RECT  197.7 204.4 198.5 215.2 ;
      RECT  195.3 205.2 196.9 206.0 ;
      RECT  196.1 204.4 196.9 205.2 ;
      RECT  190.9 225.2 191.7 214.4 ;
      RECT  194.3 215.2 195.1 214.4 ;
      RECT  196.1 223.6 196.9 214.4 ;
      RECT  192.5 225.2 193.3 214.4 ;
      RECT  197.7 225.2 198.5 214.4 ;
      RECT  195.3 224.4 196.9 223.6 ;
      RECT  196.1 225.2 196.9 224.4 ;
      RECT  190.9 225.2 191.7 236.0 ;
      RECT  194.3 235.2 195.1 236.0 ;
      RECT  196.1 226.8 196.9 236.0 ;
      RECT  192.5 225.2 193.3 236.0 ;
      RECT  197.7 225.2 198.5 236.0 ;
      RECT  195.3 226.0 196.9 226.8 ;
      RECT  196.1 225.2 196.9 226.0 ;
      RECT  190.9 246.0 191.7 235.2 ;
      RECT  194.3 236.0 195.1 235.2 ;
      RECT  196.1 244.4 196.9 235.2 ;
      RECT  192.5 246.0 193.3 235.2 ;
      RECT  197.7 246.0 198.5 235.2 ;
      RECT  195.3 245.2 196.9 244.4 ;
      RECT  196.1 246.0 196.9 245.2 ;
      RECT  190.9 246.0 191.7 256.8 ;
      RECT  194.3 256.0 195.1 256.8 ;
      RECT  196.1 247.6 196.9 256.8 ;
      RECT  192.5 246.0 193.3 256.8 ;
      RECT  197.7 246.0 198.5 256.8 ;
      RECT  195.3 246.8 196.9 247.6 ;
      RECT  196.1 246.0 196.9 246.8 ;
      RECT  190.9 266.8 191.7 256.0 ;
      RECT  194.3 256.8 195.1 256.0 ;
      RECT  196.1 265.2 196.9 256.0 ;
      RECT  192.5 266.8 193.3 256.0 ;
      RECT  197.7 266.8 198.5 256.0 ;
      RECT  195.3 266.0 196.9 265.2 ;
      RECT  196.1 266.8 196.9 266.0 ;
      RECT  190.9 266.8 191.7 277.6 ;
      RECT  194.3 276.8 195.1 277.6 ;
      RECT  196.1 268.4 196.9 277.6 ;
      RECT  192.5 266.8 193.3 277.6 ;
      RECT  197.7 266.8 198.5 277.6 ;
      RECT  195.3 267.6 196.9 268.4 ;
      RECT  196.1 266.8 196.9 267.6 ;
      RECT  190.9 287.6 191.7 276.8 ;
      RECT  194.3 277.6 195.1 276.8 ;
      RECT  196.1 286.0 196.9 276.8 ;
      RECT  192.5 287.6 193.3 276.8 ;
      RECT  197.7 287.6 198.5 276.8 ;
      RECT  195.3 286.8 196.9 286.0 ;
      RECT  196.1 287.6 196.9 286.8 ;
      RECT  190.9 287.6 191.7 298.4 ;
      RECT  194.3 297.6 195.1 298.4 ;
      RECT  196.1 289.2 196.9 298.4 ;
      RECT  192.5 287.6 193.3 298.4 ;
      RECT  197.7 287.6 198.5 298.4 ;
      RECT  195.3 288.4 196.9 289.2 ;
      RECT  196.1 287.6 196.9 288.4 ;
      RECT  190.9 308.4 191.7 297.6 ;
      RECT  194.3 298.4 195.1 297.6 ;
      RECT  196.1 306.8 196.9 297.6 ;
      RECT  192.5 308.4 193.3 297.6 ;
      RECT  197.7 308.4 198.5 297.6 ;
      RECT  195.3 307.6 196.9 306.8 ;
      RECT  196.1 308.4 196.9 307.6 ;
      RECT  190.9 308.4 191.7 319.2 ;
      RECT  194.3 318.4 195.1 319.2 ;
      RECT  196.1 310.0 196.9 319.2 ;
      RECT  192.5 308.4 193.3 319.2 ;
      RECT  197.7 308.4 198.5 319.2 ;
      RECT  195.3 309.2 196.9 310.0 ;
      RECT  196.1 308.4 196.9 309.2 ;
      RECT  190.9 329.2 191.7 318.4 ;
      RECT  194.3 319.2 195.1 318.4 ;
      RECT  196.1 327.6 196.9 318.4 ;
      RECT  192.5 329.2 193.3 318.4 ;
      RECT  197.7 329.2 198.5 318.4 ;
      RECT  195.3 328.4 196.9 327.6 ;
      RECT  196.1 329.2 196.9 328.4 ;
      RECT  190.9 329.2 191.7 340.0 ;
      RECT  194.3 339.2 195.1 340.0 ;
      RECT  196.1 330.8 196.9 340.0 ;
      RECT  192.5 329.2 193.3 340.0 ;
      RECT  197.7 329.2 198.5 340.0 ;
      RECT  195.3 330.0 196.9 330.8 ;
      RECT  196.1 329.2 196.9 330.0 ;
      RECT  190.9 350.0 191.7 339.2 ;
      RECT  194.3 340.0 195.1 339.2 ;
      RECT  196.1 348.4 196.9 339.2 ;
      RECT  192.5 350.0 193.3 339.2 ;
      RECT  197.7 350.0 198.5 339.2 ;
      RECT  195.3 349.2 196.9 348.4 ;
      RECT  196.1 350.0 196.9 349.2 ;
      RECT  185.7 183.6 186.5 350.0 ;
      RECT  189.3 183.6 190.1 350.0 ;
      RECT  192.5 183.6 193.3 350.0 ;
      RECT  196.1 183.6 196.9 350.0 ;
      RECT  187.5 297.6 188.3 298.4 ;
      RECT  187.5 297.6 188.3 298.4 ;
      RECT  194.3 276.8 195.1 277.6 ;
      RECT  194.3 297.6 195.1 298.4 ;
      RECT  187.5 193.6 188.3 194.4 ;
      RECT  194.3 297.6 195.1 298.4 ;
      RECT  187.5 339.2 188.3 340.0 ;
      RECT  194.3 193.6 195.1 194.4 ;
      RECT  194.3 318.4 195.1 319.2 ;
      RECT  194.3 318.4 195.1 319.2 ;
      RECT  194.3 339.2 195.1 340.0 ;
      RECT  194.3 235.2 195.1 236.0 ;
      RECT  194.3 235.2 195.1 236.0 ;
      RECT  187.5 214.4 188.3 215.2 ;
      RECT  187.5 276.8 188.3 277.6 ;
      RECT  187.5 235.2 188.3 236.0 ;
      RECT  187.5 235.2 188.3 236.0 ;
      RECT  187.5 256.0 188.3 256.8 ;
      RECT  194.3 256.0 195.1 256.8 ;
      RECT  187.5 318.4 188.3 319.2 ;
      RECT  187.5 318.4 188.3 319.2 ;
      RECT  194.3 214.4 195.1 215.2 ;
      RECT  184.1 214.4 184.9 225.2 ;
      RECT  197.7 256.0 198.5 266.8 ;
      RECT  190.9 276.8 191.7 287.6 ;
      RECT  190.9 276.8 191.7 287.6 ;
      RECT  197.7 339.2 198.5 350.0 ;
      RECT  184.1 339.2 184.9 350.0 ;
      RECT  190.9 266.8 191.7 277.6 ;
      RECT  190.9 266.8 191.7 277.6 ;
      RECT  190.9 225.2 191.7 236.0 ;
      RECT  190.9 225.2 191.7 236.0 ;
      RECT  197.7 266.8 198.5 277.6 ;
      RECT  197.7 287.6 198.5 298.4 ;
      RECT  197.7 214.4 198.5 225.2 ;
      RECT  190.9 308.4 191.7 319.2 ;
      RECT  190.9 308.4 191.7 319.2 ;
      RECT  184.1 204.4 184.9 215.2 ;
      RECT  184.1 193.6 184.9 204.4 ;
      RECT  184.1 225.2 184.9 236.0 ;
      RECT  190.9 214.4 191.7 225.2 ;
      RECT  190.9 214.4 191.7 225.2 ;
      RECT  197.7 297.6 198.5 308.4 ;
      RECT  190.9 256.0 191.7 266.8 ;
      RECT  190.9 256.0 191.7 266.8 ;
      RECT  184.1 266.8 184.9 277.6 ;
      RECT  197.7 308.4 198.5 319.2 ;
      RECT  197.7 204.4 198.5 215.2 ;
      RECT  184.1 235.2 184.9 246.0 ;
      RECT  184.1 297.6 184.9 308.4 ;
      RECT  184.1 246.0 184.9 256.8 ;
      RECT  184.1 318.4 184.9 329.2 ;
      RECT  190.9 204.4 191.7 215.2 ;
      RECT  190.9 204.4 191.7 215.2 ;
      RECT  184.1 183.6 184.9 194.4 ;
      RECT  190.9 193.6 191.7 204.4 ;
      RECT  190.9 193.6 191.7 204.4 ;
      RECT  190.9 246.0 191.7 256.8 ;
      RECT  190.9 183.6 191.7 194.4 ;
      RECT  197.7 235.2 198.5 246.0 ;
      RECT  190.9 246.0 191.7 256.8 ;
      RECT  184.1 308.4 184.9 319.2 ;
      RECT  184.1 329.2 184.9 340.0 ;
      RECT  190.9 287.6 191.7 298.4 ;
      RECT  190.9 287.6 191.7 298.4 ;
      RECT  190.9 318.4 191.7 329.2 ;
      RECT  190.9 318.4 191.7 329.2 ;
      RECT  184.1 276.8 184.9 287.6 ;
      RECT  197.7 225.2 198.5 236.0 ;
      RECT  190.9 339.2 191.7 350.0 ;
      RECT  190.9 339.2 191.7 350.0 ;
      RECT  197.7 276.8 198.5 287.6 ;
      RECT  190.9 297.6 191.7 308.4 ;
      RECT  190.9 297.6 191.7 308.4 ;
      RECT  190.9 329.2 191.7 340.0 ;
      RECT  190.9 329.2 191.7 340.0 ;
      RECT  197.7 318.4 198.5 329.2 ;
      RECT  190.9 235.2 191.7 246.0 ;
      RECT  190.9 235.2 191.7 246.0 ;
      RECT  184.1 256.0 184.9 266.8 ;
      RECT  197.7 183.6 198.5 194.4 ;
      RECT  197.7 193.6 198.5 204.4 ;
      RECT  197.7 246.0 198.5 256.8 ;
      RECT  184.1 287.6 184.9 298.4 ;
      RECT  197.7 329.2 198.5 340.0 ;
      RECT  190.9 183.6 191.7 194.4 ;
      RECT  184.1 162.8 184.9 173.6 ;
      RECT  177.3 162.8 178.1 173.6 ;
      RECT  180.7 172.8 181.5 173.6 ;
      RECT  182.5 162.8 183.3 173.6 ;
      RECT  178.9 162.8 179.7 173.6 ;
      RECT  177.3 183.6 178.1 172.8 ;
      RECT  180.7 173.6 181.5 172.8 ;
      RECT  182.5 182.0 183.3 172.8 ;
      RECT  178.9 183.6 179.7 172.8 ;
      RECT  184.1 183.6 184.9 172.8 ;
      RECT  181.7 182.8 183.3 182.0 ;
      RECT  182.5 183.6 183.3 182.8 ;
      RECT  177.3 183.6 178.1 194.4 ;
      RECT  180.7 193.6 181.5 194.4 ;
      RECT  182.5 185.2 183.3 194.4 ;
      RECT  178.9 183.6 179.7 194.4 ;
      RECT  184.1 183.6 184.9 194.4 ;
      RECT  181.7 184.4 183.3 185.2 ;
      RECT  182.5 183.6 183.3 184.4 ;
      RECT  177.3 204.4 178.1 193.6 ;
      RECT  180.7 194.4 181.5 193.6 ;
      RECT  182.5 202.8 183.3 193.6 ;
      RECT  178.9 204.4 179.7 193.6 ;
      RECT  184.1 204.4 184.9 193.6 ;
      RECT  181.7 203.6 183.3 202.8 ;
      RECT  182.5 204.4 183.3 203.6 ;
      RECT  177.3 204.4 178.1 215.2 ;
      RECT  180.7 214.4 181.5 215.2 ;
      RECT  182.5 206.0 183.3 215.2 ;
      RECT  178.9 204.4 179.7 215.2 ;
      RECT  184.1 204.4 184.9 215.2 ;
      RECT  181.7 205.2 183.3 206.0 ;
      RECT  182.5 204.4 183.3 205.2 ;
      RECT  177.3 225.2 178.1 214.4 ;
      RECT  180.7 215.2 181.5 214.4 ;
      RECT  182.5 223.6 183.3 214.4 ;
      RECT  178.9 225.2 179.7 214.4 ;
      RECT  184.1 225.2 184.9 214.4 ;
      RECT  181.7 224.4 183.3 223.6 ;
      RECT  182.5 225.2 183.3 224.4 ;
      RECT  177.3 225.2 178.1 236.0 ;
      RECT  180.7 235.2 181.5 236.0 ;
      RECT  182.5 226.8 183.3 236.0 ;
      RECT  178.9 225.2 179.7 236.0 ;
      RECT  184.1 225.2 184.9 236.0 ;
      RECT  181.7 226.0 183.3 226.8 ;
      RECT  182.5 225.2 183.3 226.0 ;
      RECT  177.3 246.0 178.1 235.2 ;
      RECT  180.7 236.0 181.5 235.2 ;
      RECT  182.5 244.4 183.3 235.2 ;
      RECT  178.9 246.0 179.7 235.2 ;
      RECT  184.1 246.0 184.9 235.2 ;
      RECT  181.7 245.2 183.3 244.4 ;
      RECT  182.5 246.0 183.3 245.2 ;
      RECT  177.3 246.0 178.1 256.8 ;
      RECT  180.7 256.0 181.5 256.8 ;
      RECT  182.5 247.6 183.3 256.8 ;
      RECT  178.9 246.0 179.7 256.8 ;
      RECT  184.1 246.0 184.9 256.8 ;
      RECT  181.7 246.8 183.3 247.6 ;
      RECT  182.5 246.0 183.3 246.8 ;
      RECT  177.3 266.8 178.1 256.0 ;
      RECT  180.7 256.8 181.5 256.0 ;
      RECT  182.5 265.2 183.3 256.0 ;
      RECT  178.9 266.8 179.7 256.0 ;
      RECT  184.1 266.8 184.9 256.0 ;
      RECT  181.7 266.0 183.3 265.2 ;
      RECT  182.5 266.8 183.3 266.0 ;
      RECT  177.3 266.8 178.1 277.6 ;
      RECT  180.7 276.8 181.5 277.6 ;
      RECT  182.5 268.4 183.3 277.6 ;
      RECT  178.9 266.8 179.7 277.6 ;
      RECT  184.1 266.8 184.9 277.6 ;
      RECT  181.7 267.6 183.3 268.4 ;
      RECT  182.5 266.8 183.3 267.6 ;
      RECT  177.3 287.6 178.1 276.8 ;
      RECT  180.7 277.6 181.5 276.8 ;
      RECT  182.5 286.0 183.3 276.8 ;
      RECT  178.9 287.6 179.7 276.8 ;
      RECT  184.1 287.6 184.9 276.8 ;
      RECT  181.7 286.8 183.3 286.0 ;
      RECT  182.5 287.6 183.3 286.8 ;
      RECT  177.3 287.6 178.1 298.4 ;
      RECT  180.7 297.6 181.5 298.4 ;
      RECT  182.5 289.2 183.3 298.4 ;
      RECT  178.9 287.6 179.7 298.4 ;
      RECT  184.1 287.6 184.9 298.4 ;
      RECT  181.7 288.4 183.3 289.2 ;
      RECT  182.5 287.6 183.3 288.4 ;
      RECT  177.3 308.4 178.1 297.6 ;
      RECT  180.7 298.4 181.5 297.6 ;
      RECT  182.5 306.8 183.3 297.6 ;
      RECT  178.9 308.4 179.7 297.6 ;
      RECT  184.1 308.4 184.9 297.6 ;
      RECT  181.7 307.6 183.3 306.8 ;
      RECT  182.5 308.4 183.3 307.6 ;
      RECT  177.3 308.4 178.1 319.2 ;
      RECT  180.7 318.4 181.5 319.2 ;
      RECT  182.5 310.0 183.3 319.2 ;
      RECT  178.9 308.4 179.7 319.2 ;
      RECT  184.1 308.4 184.9 319.2 ;
      RECT  181.7 309.2 183.3 310.0 ;
      RECT  182.5 308.4 183.3 309.2 ;
      RECT  177.3 329.2 178.1 318.4 ;
      RECT  180.7 319.2 181.5 318.4 ;
      RECT  182.5 327.6 183.3 318.4 ;
      RECT  178.9 329.2 179.7 318.4 ;
      RECT  184.1 329.2 184.9 318.4 ;
      RECT  181.7 328.4 183.3 327.6 ;
      RECT  182.5 329.2 183.3 328.4 ;
      RECT  177.3 329.2 178.1 340.0 ;
      RECT  180.7 339.2 181.5 340.0 ;
      RECT  182.5 330.8 183.3 340.0 ;
      RECT  178.9 329.2 179.7 340.0 ;
      RECT  184.1 329.2 184.9 340.0 ;
      RECT  181.7 330.0 183.3 330.8 ;
      RECT  182.5 329.2 183.3 330.0 ;
      RECT  177.3 350.0 178.1 339.2 ;
      RECT  180.7 340.0 181.5 339.2 ;
      RECT  182.5 348.4 183.3 339.2 ;
      RECT  178.9 350.0 179.7 339.2 ;
      RECT  184.1 350.0 184.9 339.2 ;
      RECT  181.7 349.2 183.3 348.4 ;
      RECT  182.5 350.0 183.3 349.2 ;
      RECT  184.1 350.0 184.9 360.8 ;
      RECT  177.3 350.0 178.1 360.8 ;
      RECT  180.7 360.0 181.5 360.8 ;
      RECT  182.5 350.0 183.3 360.8 ;
      RECT  178.9 350.0 179.7 360.8 ;
      RECT  180.7 214.4 181.5 215.2 ;
      RECT  180.7 214.4 181.5 215.2 ;
      RECT  180.7 339.2 181.5 340.0 ;
      RECT  180.7 276.8 181.5 277.6 ;
      RECT  180.7 276.8 181.5 277.6 ;
      RECT  180.7 297.6 181.5 298.4 ;
      RECT  180.7 172.8 181.5 173.6 ;
      RECT  180.7 235.2 181.5 236.0 ;
      RECT  180.7 193.6 181.5 194.4 ;
      RECT  180.7 318.4 181.5 319.2 ;
      RECT  180.7 297.6 181.5 298.4 ;
      RECT  180.7 256.0 181.5 256.8 ;
      RECT  177.3 193.6 178.1 204.4 ;
      RECT  184.1 256.0 184.9 266.8 ;
      RECT  177.3 318.4 178.1 329.2 ;
      RECT  184.1 246.0 184.9 256.8 ;
      RECT  184.1 204.4 184.9 215.2 ;
      RECT  184.1 287.6 184.9 298.4 ;
      RECT  184.1 329.2 184.9 340.0 ;
      RECT  177.3 183.6 178.1 194.4 ;
      RECT  177.3 172.8 178.1 183.6 ;
      RECT  177.3 204.4 178.1 215.2 ;
      RECT  184.1 193.6 184.9 204.4 ;
      RECT  184.1 235.2 184.9 246.0 ;
      RECT  177.3 246.0 178.1 256.8 ;
      RECT  177.3 214.4 178.1 225.2 ;
      RECT  177.3 276.8 178.1 287.6 ;
      RECT  177.3 225.2 178.1 236.0 ;
      RECT  177.3 297.6 178.1 308.4 ;
      RECT  184.1 183.6 184.9 194.4 ;
      RECT  184.1 172.8 184.9 183.6 ;
      RECT  177.3 308.4 178.1 319.2 ;
      RECT  184.1 225.2 184.9 236.0 ;
      RECT  177.3 287.6 178.1 298.4 ;
      RECT  184.1 266.8 184.9 277.6 ;
      RECT  184.1 297.6 184.9 308.4 ;
      RECT  177.3 256.0 178.1 266.8 ;
      RECT  184.1 318.4 184.9 329.2 ;
      RECT  184.1 308.4 184.9 319.2 ;
      RECT  184.1 276.8 184.9 287.6 ;
      RECT  177.3 329.2 178.1 340.0 ;
      RECT  184.1 214.4 184.9 225.2 ;
      RECT  177.3 235.2 178.1 246.0 ;
      RECT  177.3 339.2 178.1 350.0 ;
      RECT  184.1 339.2 184.9 350.0 ;
      RECT  177.3 266.8 178.1 277.6 ;
      RECT  190.9 183.6 191.7 172.8 ;
      RECT  184.1 183.6 184.9 172.8 ;
      RECT  187.5 173.6 188.3 172.8 ;
      RECT  189.3 183.6 190.1 172.8 ;
      RECT  185.7 183.6 186.5 172.8 ;
      RECT  197.7 183.6 198.5 172.8 ;
      RECT  190.9 183.6 191.7 172.8 ;
      RECT  194.3 173.6 195.1 172.8 ;
      RECT  196.1 183.6 196.9 172.8 ;
      RECT  192.5 183.6 193.3 172.8 ;
      RECT  185.7 183.6 186.5 173.2 ;
      RECT  189.3 183.6 190.1 173.2 ;
      RECT  192.5 183.6 193.3 173.2 ;
      RECT  196.1 183.6 196.9 173.2 ;
      RECT  187.5 173.6 188.3 172.8 ;
      RECT  194.3 173.6 195.1 172.8 ;
      RECT  197.7 183.6 198.5 172.8 ;
      RECT  184.1 183.6 184.9 172.8 ;
      RECT  190.9 183.6 191.7 172.8 ;
      RECT  190.9 183.6 191.7 172.8 ;
      RECT  190.9 162.8 191.7 173.6 ;
      RECT  184.1 162.8 184.9 173.6 ;
      RECT  187.5 172.8 188.3 173.6 ;
      RECT  189.3 162.8 190.1 173.6 ;
      RECT  185.7 162.8 186.5 173.6 ;
      RECT  197.7 162.8 198.5 173.6 ;
      RECT  190.9 162.8 191.7 173.6 ;
      RECT  194.3 172.8 195.1 173.6 ;
      RECT  196.1 162.8 196.9 173.6 ;
      RECT  192.5 162.8 193.3 173.6 ;
      RECT  185.7 162.8 186.5 173.2 ;
      RECT  189.3 162.8 190.1 173.2 ;
      RECT  192.5 162.8 193.3 173.2 ;
      RECT  196.1 162.8 196.9 173.2 ;
      RECT  187.5 172.8 188.3 173.6 ;
      RECT  194.3 172.8 195.1 173.6 ;
      RECT  197.7 162.8 198.5 173.6 ;
      RECT  184.1 162.8 184.9 173.6 ;
      RECT  190.9 162.8 191.7 173.6 ;
      RECT  190.9 162.8 191.7 173.6 ;
      RECT  190.9 350.0 191.7 360.8 ;
      RECT  184.1 350.0 184.9 360.8 ;
      RECT  187.5 360.0 188.3 360.8 ;
      RECT  189.3 350.0 190.1 360.8 ;
      RECT  185.7 350.0 186.5 360.8 ;
      RECT  197.7 350.0 198.5 360.8 ;
      RECT  190.9 350.0 191.7 360.8 ;
      RECT  194.3 360.0 195.1 360.8 ;
      RECT  196.1 350.0 196.9 360.8 ;
      RECT  192.5 350.0 193.3 360.8 ;
      RECT  185.7 350.0 186.5 360.4 ;
      RECT  189.3 350.0 190.1 360.4 ;
      RECT  192.5 350.0 193.3 360.4 ;
      RECT  196.1 350.0 196.9 360.4 ;
      RECT  187.5 360.0 188.3 360.8 ;
      RECT  194.3 360.0 195.1 360.8 ;
      RECT  197.7 350.0 198.5 360.8 ;
      RECT  184.1 350.0 184.9 360.8 ;
      RECT  190.9 350.0 191.7 360.8 ;
      RECT  190.9 350.0 191.7 360.8 ;
      RECT  177.3 162.8 178.1 173.6 ;
      RECT  170.5 162.8 171.3 173.6 ;
      RECT  173.9 172.8 174.7 173.6 ;
      RECT  175.7 162.8 176.5 173.6 ;
      RECT  172.1 162.8 172.9 173.6 ;
      RECT  177.3 183.6 178.1 172.8 ;
      RECT  170.5 183.6 171.3 172.8 ;
      RECT  173.9 173.6 174.7 172.8 ;
      RECT  175.7 183.6 176.5 172.8 ;
      RECT  172.1 183.6 172.9 172.8 ;
      RECT  177.3 183.6 178.1 194.4 ;
      RECT  170.5 183.6 171.3 194.4 ;
      RECT  173.9 193.6 174.7 194.4 ;
      RECT  175.7 183.6 176.5 194.4 ;
      RECT  172.1 183.6 172.9 194.4 ;
      RECT  177.3 204.4 178.1 193.6 ;
      RECT  170.5 204.4 171.3 193.6 ;
      RECT  173.9 194.4 174.7 193.6 ;
      RECT  175.7 204.4 176.5 193.6 ;
      RECT  172.1 204.4 172.9 193.6 ;
      RECT  177.3 204.4 178.1 215.2 ;
      RECT  170.5 204.4 171.3 215.2 ;
      RECT  173.9 214.4 174.7 215.2 ;
      RECT  175.7 204.4 176.5 215.2 ;
      RECT  172.1 204.4 172.9 215.2 ;
      RECT  177.3 225.2 178.1 214.4 ;
      RECT  170.5 225.2 171.3 214.4 ;
      RECT  173.9 215.2 174.7 214.4 ;
      RECT  175.7 225.2 176.5 214.4 ;
      RECT  172.1 225.2 172.9 214.4 ;
      RECT  177.3 225.2 178.1 236.0 ;
      RECT  170.5 225.2 171.3 236.0 ;
      RECT  173.9 235.2 174.7 236.0 ;
      RECT  175.7 225.2 176.5 236.0 ;
      RECT  172.1 225.2 172.9 236.0 ;
      RECT  177.3 246.0 178.1 235.2 ;
      RECT  170.5 246.0 171.3 235.2 ;
      RECT  173.9 236.0 174.7 235.2 ;
      RECT  175.7 246.0 176.5 235.2 ;
      RECT  172.1 246.0 172.9 235.2 ;
      RECT  177.3 246.0 178.1 256.8 ;
      RECT  170.5 246.0 171.3 256.8 ;
      RECT  173.9 256.0 174.7 256.8 ;
      RECT  175.7 246.0 176.5 256.8 ;
      RECT  172.1 246.0 172.9 256.8 ;
      RECT  177.3 266.8 178.1 256.0 ;
      RECT  170.5 266.8 171.3 256.0 ;
      RECT  173.9 256.8 174.7 256.0 ;
      RECT  175.7 266.8 176.5 256.0 ;
      RECT  172.1 266.8 172.9 256.0 ;
      RECT  177.3 266.8 178.1 277.6 ;
      RECT  170.5 266.8 171.3 277.6 ;
      RECT  173.9 276.8 174.7 277.6 ;
      RECT  175.7 266.8 176.5 277.6 ;
      RECT  172.1 266.8 172.9 277.6 ;
      RECT  177.3 287.6 178.1 276.8 ;
      RECT  170.5 287.6 171.3 276.8 ;
      RECT  173.9 277.6 174.7 276.8 ;
      RECT  175.7 287.6 176.5 276.8 ;
      RECT  172.1 287.6 172.9 276.8 ;
      RECT  177.3 287.6 178.1 298.4 ;
      RECT  170.5 287.6 171.3 298.4 ;
      RECT  173.9 297.6 174.7 298.4 ;
      RECT  175.7 287.6 176.5 298.4 ;
      RECT  172.1 287.6 172.9 298.4 ;
      RECT  177.3 308.4 178.1 297.6 ;
      RECT  170.5 308.4 171.3 297.6 ;
      RECT  173.9 298.4 174.7 297.6 ;
      RECT  175.7 308.4 176.5 297.6 ;
      RECT  172.1 308.4 172.9 297.6 ;
      RECT  177.3 308.4 178.1 319.2 ;
      RECT  170.5 308.4 171.3 319.2 ;
      RECT  173.9 318.4 174.7 319.2 ;
      RECT  175.7 308.4 176.5 319.2 ;
      RECT  172.1 308.4 172.9 319.2 ;
      RECT  177.3 329.2 178.1 318.4 ;
      RECT  170.5 329.2 171.3 318.4 ;
      RECT  173.9 319.2 174.7 318.4 ;
      RECT  175.7 329.2 176.5 318.4 ;
      RECT  172.1 329.2 172.9 318.4 ;
      RECT  177.3 329.2 178.1 340.0 ;
      RECT  170.5 329.2 171.3 340.0 ;
      RECT  173.9 339.2 174.7 340.0 ;
      RECT  175.7 329.2 176.5 340.0 ;
      RECT  172.1 329.2 172.9 340.0 ;
      RECT  177.3 350.0 178.1 339.2 ;
      RECT  170.5 350.0 171.3 339.2 ;
      RECT  173.9 340.0 174.7 339.2 ;
      RECT  175.7 350.0 176.5 339.2 ;
      RECT  172.1 350.0 172.9 339.2 ;
      RECT  177.3 350.0 178.1 360.8 ;
      RECT  170.5 350.0 171.3 360.8 ;
      RECT  173.9 360.0 174.7 360.8 ;
      RECT  175.7 350.0 176.5 360.8 ;
      RECT  172.1 350.0 172.9 360.8 ;
      RECT  172.1 162.8 172.9 360.4 ;
      RECT  175.7 162.8 176.5 360.4 ;
      RECT  173.9 214.4 174.7 215.2 ;
      RECT  173.9 214.4 174.7 215.2 ;
      RECT  173.9 339.2 174.7 340.0 ;
      RECT  173.9 360.0 174.7 360.8 ;
      RECT  173.9 276.8 174.7 277.6 ;
      RECT  173.9 276.8 174.7 277.6 ;
      RECT  173.9 297.6 174.7 298.4 ;
      RECT  173.9 172.8 174.7 173.6 ;
      RECT  173.9 235.2 174.7 236.0 ;
      RECT  173.9 193.6 174.7 194.4 ;
      RECT  173.9 318.4 174.7 319.2 ;
      RECT  173.9 297.6 174.7 298.4 ;
      RECT  173.9 256.0 174.7 256.8 ;
      RECT  170.5 193.6 171.3 204.4 ;
      RECT  177.3 256.0 178.1 266.8 ;
      RECT  170.5 318.4 171.3 329.2 ;
      RECT  177.3 246.0 178.1 256.8 ;
      RECT  177.3 204.4 178.1 215.2 ;
      RECT  177.3 287.6 178.1 298.4 ;
      RECT  177.3 350.0 178.1 360.8 ;
      RECT  177.3 329.2 178.1 340.0 ;
      RECT  170.5 183.6 171.3 194.4 ;
      RECT  170.5 172.8 171.3 183.6 ;
      RECT  170.5 204.4 171.3 215.2 ;
      RECT  177.3 193.6 178.1 204.4 ;
      RECT  177.3 235.2 178.1 246.0 ;
      RECT  170.5 246.0 171.3 256.8 ;
      RECT  170.5 214.4 171.3 225.2 ;
      RECT  170.5 276.8 171.3 287.6 ;
      RECT  170.5 225.2 171.3 236.0 ;
      RECT  170.5 297.6 171.3 308.4 ;
      RECT  177.3 183.6 178.1 194.4 ;
      RECT  170.5 162.8 171.3 173.6 ;
      RECT  177.3 172.8 178.1 183.6 ;
      RECT  170.5 308.4 171.3 319.2 ;
      RECT  177.3 225.2 178.1 236.0 ;
      RECT  170.5 287.6 171.3 298.4 ;
      RECT  170.5 350.0 171.3 360.8 ;
      RECT  177.3 266.8 178.1 277.6 ;
      RECT  177.3 297.6 178.1 308.4 ;
      RECT  170.5 256.0 171.3 266.8 ;
      RECT  177.3 318.4 178.1 329.2 ;
      RECT  177.3 308.4 178.1 319.2 ;
      RECT  177.3 276.8 178.1 287.6 ;
      RECT  170.5 329.2 171.3 340.0 ;
      RECT  177.3 214.4 178.1 225.2 ;
      RECT  170.5 235.2 171.3 246.0 ;
      RECT  170.5 339.2 171.3 350.0 ;
      RECT  177.3 339.2 178.1 350.0 ;
      RECT  170.5 266.8 171.3 277.6 ;
      RECT  177.3 162.8 178.1 173.6 ;
      RECT  204.5 162.8 205.3 173.6 ;
      RECT  197.7 162.8 198.5 173.6 ;
      RECT  201.1 172.8 201.9 173.6 ;
      RECT  202.9 162.8 203.7 173.6 ;
      RECT  199.3 162.8 200.1 173.6 ;
      RECT  204.5 183.6 205.3 172.8 ;
      RECT  197.7 183.6 198.5 172.8 ;
      RECT  201.1 173.6 201.9 172.8 ;
      RECT  202.9 183.6 203.7 172.8 ;
      RECT  199.3 183.6 200.1 172.8 ;
      RECT  204.5 183.6 205.3 194.4 ;
      RECT  197.7 183.6 198.5 194.4 ;
      RECT  201.1 193.6 201.9 194.4 ;
      RECT  202.9 183.6 203.7 194.4 ;
      RECT  199.3 183.6 200.1 194.4 ;
      RECT  204.5 204.4 205.3 193.6 ;
      RECT  197.7 204.4 198.5 193.6 ;
      RECT  201.1 194.4 201.9 193.6 ;
      RECT  202.9 204.4 203.7 193.6 ;
      RECT  199.3 204.4 200.1 193.6 ;
      RECT  204.5 204.4 205.3 215.2 ;
      RECT  197.7 204.4 198.5 215.2 ;
      RECT  201.1 214.4 201.9 215.2 ;
      RECT  202.9 204.4 203.7 215.2 ;
      RECT  199.3 204.4 200.1 215.2 ;
      RECT  204.5 225.2 205.3 214.4 ;
      RECT  197.7 225.2 198.5 214.4 ;
      RECT  201.1 215.2 201.9 214.4 ;
      RECT  202.9 225.2 203.7 214.4 ;
      RECT  199.3 225.2 200.1 214.4 ;
      RECT  204.5 225.2 205.3 236.0 ;
      RECT  197.7 225.2 198.5 236.0 ;
      RECT  201.1 235.2 201.9 236.0 ;
      RECT  202.9 225.2 203.7 236.0 ;
      RECT  199.3 225.2 200.1 236.0 ;
      RECT  204.5 246.0 205.3 235.2 ;
      RECT  197.7 246.0 198.5 235.2 ;
      RECT  201.1 236.0 201.9 235.2 ;
      RECT  202.9 246.0 203.7 235.2 ;
      RECT  199.3 246.0 200.1 235.2 ;
      RECT  204.5 246.0 205.3 256.8 ;
      RECT  197.7 246.0 198.5 256.8 ;
      RECT  201.1 256.0 201.9 256.8 ;
      RECT  202.9 246.0 203.7 256.8 ;
      RECT  199.3 246.0 200.1 256.8 ;
      RECT  204.5 266.8 205.3 256.0 ;
      RECT  197.7 266.8 198.5 256.0 ;
      RECT  201.1 256.8 201.9 256.0 ;
      RECT  202.9 266.8 203.7 256.0 ;
      RECT  199.3 266.8 200.1 256.0 ;
      RECT  204.5 266.8 205.3 277.6 ;
      RECT  197.7 266.8 198.5 277.6 ;
      RECT  201.1 276.8 201.9 277.6 ;
      RECT  202.9 266.8 203.7 277.6 ;
      RECT  199.3 266.8 200.1 277.6 ;
      RECT  204.5 287.6 205.3 276.8 ;
      RECT  197.7 287.6 198.5 276.8 ;
      RECT  201.1 277.6 201.9 276.8 ;
      RECT  202.9 287.6 203.7 276.8 ;
      RECT  199.3 287.6 200.1 276.8 ;
      RECT  204.5 287.6 205.3 298.4 ;
      RECT  197.7 287.6 198.5 298.4 ;
      RECT  201.1 297.6 201.9 298.4 ;
      RECT  202.9 287.6 203.7 298.4 ;
      RECT  199.3 287.6 200.1 298.4 ;
      RECT  204.5 308.4 205.3 297.6 ;
      RECT  197.7 308.4 198.5 297.6 ;
      RECT  201.1 298.4 201.9 297.6 ;
      RECT  202.9 308.4 203.7 297.6 ;
      RECT  199.3 308.4 200.1 297.6 ;
      RECT  204.5 308.4 205.3 319.2 ;
      RECT  197.7 308.4 198.5 319.2 ;
      RECT  201.1 318.4 201.9 319.2 ;
      RECT  202.9 308.4 203.7 319.2 ;
      RECT  199.3 308.4 200.1 319.2 ;
      RECT  204.5 329.2 205.3 318.4 ;
      RECT  197.7 329.2 198.5 318.4 ;
      RECT  201.1 319.2 201.9 318.4 ;
      RECT  202.9 329.2 203.7 318.4 ;
      RECT  199.3 329.2 200.1 318.4 ;
      RECT  204.5 329.2 205.3 340.0 ;
      RECT  197.7 329.2 198.5 340.0 ;
      RECT  201.1 339.2 201.9 340.0 ;
      RECT  202.9 329.2 203.7 340.0 ;
      RECT  199.3 329.2 200.1 340.0 ;
      RECT  204.5 350.0 205.3 339.2 ;
      RECT  197.7 350.0 198.5 339.2 ;
      RECT  201.1 340.0 201.9 339.2 ;
      RECT  202.9 350.0 203.7 339.2 ;
      RECT  199.3 350.0 200.1 339.2 ;
      RECT  204.5 350.0 205.3 360.8 ;
      RECT  197.7 350.0 198.5 360.8 ;
      RECT  201.1 360.0 201.9 360.8 ;
      RECT  202.9 350.0 203.7 360.8 ;
      RECT  199.3 350.0 200.1 360.8 ;
      RECT  199.3 162.8 200.1 360.4 ;
      RECT  202.9 162.8 203.7 360.4 ;
      RECT  201.1 214.4 201.9 215.2 ;
      RECT  201.1 214.4 201.9 215.2 ;
      RECT  201.1 339.2 201.9 340.0 ;
      RECT  201.1 360.0 201.9 360.8 ;
      RECT  201.1 276.8 201.9 277.6 ;
      RECT  201.1 276.8 201.9 277.6 ;
      RECT  201.1 297.6 201.9 298.4 ;
      RECT  201.1 172.8 201.9 173.6 ;
      RECT  201.1 235.2 201.9 236.0 ;
      RECT  201.1 193.6 201.9 194.4 ;
      RECT  201.1 318.4 201.9 319.2 ;
      RECT  201.1 297.6 201.9 298.4 ;
      RECT  201.1 256.0 201.9 256.8 ;
      RECT  197.7 193.6 198.5 204.4 ;
      RECT  204.5 256.0 205.3 266.8 ;
      RECT  197.7 318.4 198.5 329.2 ;
      RECT  204.5 246.0 205.3 256.8 ;
      RECT  204.5 204.4 205.3 215.2 ;
      RECT  204.5 287.6 205.3 298.4 ;
      RECT  204.5 350.0 205.3 360.8 ;
      RECT  204.5 329.2 205.3 340.0 ;
      RECT  197.7 183.6 198.5 194.4 ;
      RECT  197.7 172.8 198.5 183.6 ;
      RECT  197.7 204.4 198.5 215.2 ;
      RECT  204.5 193.6 205.3 204.4 ;
      RECT  204.5 235.2 205.3 246.0 ;
      RECT  197.7 246.0 198.5 256.8 ;
      RECT  197.7 214.4 198.5 225.2 ;
      RECT  197.7 276.8 198.5 287.6 ;
      RECT  197.7 225.2 198.5 236.0 ;
      RECT  197.7 297.6 198.5 308.4 ;
      RECT  204.5 183.6 205.3 194.4 ;
      RECT  197.7 162.8 198.5 173.6 ;
      RECT  204.5 172.8 205.3 183.6 ;
      RECT  197.7 308.4 198.5 319.2 ;
      RECT  204.5 225.2 205.3 236.0 ;
      RECT  197.7 287.6 198.5 298.4 ;
      RECT  197.7 350.0 198.5 360.8 ;
      RECT  204.5 266.8 205.3 277.6 ;
      RECT  204.5 297.6 205.3 308.4 ;
      RECT  197.7 256.0 198.5 266.8 ;
      RECT  204.5 318.4 205.3 329.2 ;
      RECT  204.5 308.4 205.3 319.2 ;
      RECT  204.5 276.8 205.3 287.6 ;
      RECT  197.7 329.2 198.5 340.0 ;
      RECT  204.5 214.4 205.3 225.2 ;
      RECT  197.7 235.2 198.5 246.0 ;
      RECT  197.7 339.2 198.5 350.0 ;
      RECT  204.5 339.2 205.3 350.0 ;
      RECT  197.7 266.8 198.5 277.6 ;
      RECT  204.5 162.8 205.3 173.6 ;
      RECT  185.7 162.8 186.5 360.4 ;
      RECT  189.3 162.8 190.1 360.4 ;
      RECT  192.5 162.8 193.3 360.4 ;
      RECT  196.1 162.8 196.9 360.4 ;
      RECT  178.9 162.8 179.7 360.4 ;
      RECT  182.5 162.8 183.3 360.4 ;
      RECT  180.7 256.0 181.5 256.8 ;
      RECT  180.7 276.8 181.5 277.6 ;
      RECT  180.7 339.2 181.5 340.0 ;
      RECT  180.7 172.8 181.5 173.6 ;
      RECT  180.7 297.6 181.5 298.4 ;
      RECT  180.7 318.4 181.5 319.2 ;
      RECT  180.7 214.4 181.5 215.2 ;
      RECT  180.7 235.2 181.5 236.0 ;
      RECT  180.7 193.6 181.5 194.4 ;
      RECT  184.1 235.2 184.9 246.0 ;
      RECT  177.3 256.0 178.1 266.8 ;
      RECT  184.1 318.4 184.9 329.2 ;
      RECT  184.1 246.0 184.9 256.8 ;
      RECT  177.3 193.6 178.1 204.4 ;
      RECT  177.3 235.2 178.1 246.0 ;
      RECT  177.3 183.6 178.1 194.4 ;
      RECT  177.3 297.6 178.1 308.4 ;
      RECT  177.3 318.4 178.1 329.2 ;
      RECT  177.3 276.8 178.1 287.6 ;
      RECT  184.1 297.6 184.9 308.4 ;
      RECT  177.3 287.6 178.1 298.4 ;
      RECT  184.1 276.8 184.9 287.6 ;
      RECT  177.3 172.8 178.1 183.6 ;
      RECT  184.1 308.4 184.9 319.2 ;
      RECT  177.3 246.0 178.1 256.8 ;
      RECT  177.3 204.4 178.1 215.2 ;
      RECT  184.1 266.8 184.9 277.6 ;
      RECT  184.1 193.6 184.9 204.4 ;
      RECT  184.1 287.6 184.9 298.4 ;
      RECT  184.1 329.2 184.9 340.0 ;
      RECT  177.3 225.2 178.1 236.0 ;
      RECT  184.1 204.4 184.9 215.2 ;
      RECT  184.1 256.0 184.9 266.8 ;
      RECT  177.3 308.4 178.1 319.2 ;
      RECT  184.1 225.2 184.9 236.0 ;
      RECT  177.3 329.2 178.1 340.0 ;
      RECT  184.1 183.6 184.9 194.4 ;
      RECT  184.1 214.4 184.9 225.2 ;
      RECT  177.3 266.8 178.1 277.6 ;
      RECT  184.1 339.2 184.9 350.0 ;
      RECT  177.3 214.4 178.1 225.2 ;
      RECT  184.1 172.8 184.9 183.6 ;
      RECT  177.3 339.2 178.1 350.0 ;
      RECT  178.8 146.6 179.4 158.6 ;
      RECT  182.8 146.6 183.4 158.6 ;
      RECT  185.6 146.6 186.2 158.6 ;
      RECT  189.6 146.6 190.2 158.6 ;
      RECT  192.4 146.6 193.0 158.6 ;
      RECT  196.4 146.6 197.0 158.6 ;
      RECT  178.8 146.6 179.4 158.6 ;
      RECT  182.8 146.6 183.4 158.6 ;
      RECT  185.6 146.6 186.2 158.6 ;
      RECT  189.6 146.6 190.2 158.6 ;
      RECT  192.4 146.6 193.0 158.6 ;
      RECT  196.4 146.6 197.0 158.6 ;
      RECT  189.9 122.2 190.7 123.8 ;
      RECT  188.5 118.6 189.7 119.4 ;
      RECT  186.5 118.6 187.9 119.4 ;
      RECT  186.5 119.4 187.3 142.4 ;
      RECT  188.5 119.4 189.3 142.4 ;
      RECT  190.9 135.6 191.7 137.2 ;
      RECT  186.5 109.8 187.3 118.6 ;
      RECT  188.5 109.8 189.3 118.6 ;
      RECT  185.1 109.8 185.9 112.8 ;
      RECT  196.7 122.2 197.5 123.8 ;
      RECT  195.3 118.6 196.5 119.4 ;
      RECT  193.3 118.6 194.7 119.4 ;
      RECT  193.3 119.4 194.1 142.4 ;
      RECT  195.3 119.4 196.1 142.4 ;
      RECT  197.7 135.6 198.5 137.2 ;
      RECT  193.3 109.8 194.1 118.6 ;
      RECT  195.3 109.8 196.1 118.6 ;
      RECT  191.9 109.8 192.7 112.8 ;
      RECT  185.1 109.8 185.9 112.8 ;
      RECT  186.5 119.4 187.3 142.4 ;
      RECT  188.5 119.4 189.3 142.4 ;
      RECT  191.9 109.8 192.7 112.8 ;
      RECT  193.3 119.4 194.1 142.4 ;
      RECT  195.3 119.4 196.1 142.4 ;
      RECT  186.5 103.6 187.3 105.6 ;
      RECT  188.3 77.8 189.1 78.6 ;
      RECT  188.3 71.2 189.1 72.0 ;
      RECT  186.9 96.8 187.7 97.6 ;
      RECT  189.7 82.2 190.5 83.0 ;
      RECT  187.7 88.6 188.5 89.4 ;
      RECT  187.5 65.0 188.3 67.0 ;
      RECT  188.5 100.6 189.3 105.6 ;
      RECT  193.3 103.6 194.1 105.6 ;
      RECT  195.1 77.8 195.9 78.6 ;
      RECT  195.1 71.2 195.9 72.0 ;
      RECT  193.7 96.8 194.5 97.6 ;
      RECT  196.5 82.2 197.3 83.0 ;
      RECT  194.5 88.6 195.3 89.4 ;
      RECT  194.3 65.0 195.1 67.0 ;
      RECT  195.3 100.6 196.1 105.6 ;
      RECT  187.5 65.0 188.3 67.0 ;
      RECT  194.3 65.0 195.1 67.0 ;
      RECT  186.5 103.6 187.3 105.6 ;
      RECT  188.5 100.6 189.3 105.6 ;
      RECT  193.3 103.6 194.1 105.6 ;
      RECT  195.3 100.6 196.1 105.6 ;
      RECT  178.8 158.6 179.4 146.6 ;
      RECT  182.8 158.6 183.4 146.6 ;
      RECT  185.6 158.6 186.2 146.6 ;
      RECT  189.6 158.6 190.2 146.6 ;
      RECT  192.4 158.6 193.0 146.6 ;
      RECT  196.4 158.6 197.0 146.6 ;
      RECT  185.1 112.8 185.9 109.8 ;
      RECT  191.9 112.8 192.7 109.8 ;
      RECT  187.5 67.0 188.3 65.0 ;
      RECT  194.3 67.0 195.1 65.0 ;
      RECT  87.4 188.6 88.2 189.4 ;
      RECT  88.8 199.4 89.6 200.2 ;
      RECT  87.4 251.0 88.2 251.8 ;
      RECT  88.8 261.8 89.6 262.6 ;
      RECT  79.9 184.0 80.5 288.0 ;
      RECT  81.3 184.0 81.9 288.0 ;
      RECT  82.7 184.0 83.3 288.0 ;
      RECT  84.1 184.0 84.7 288.0 ;
      RECT  154.5 184.0 155.1 350.4 ;
      RECT  79.9 184.0 80.5 288.0 ;
      RECT  81.3 184.0 81.9 288.0 ;
      RECT  82.7 184.0 83.3 288.0 ;
      RECT  84.1 184.0 84.7 288.0 ;
      RECT  154.5 184.0 155.1 350.4 ;
      RECT  185.1 109.8 185.9 112.8 ;
      RECT  191.9 109.8 192.7 112.8 ;
      RECT  187.5 65.0 188.3 67.0 ;
      RECT  194.3 65.0 195.1 67.0 ;
      RECT  79.9 184.0 80.5 288.0 ;
      RECT  81.3 184.0 81.9 288.0 ;
      RECT  82.7 184.0 83.3 288.0 ;
      RECT  84.1 184.0 84.7 288.0 ;
      RECT  163.9 65.0 164.5 180.8 ;
      RECT  166.7 65.0 167.3 180.8 ;
      RECT  165.3 65.0 165.9 180.8 ;
      RECT  168.1 65.0 168.7 180.8 ;
      RECT  4.4 3.2 5.2 14.8 ;
      RECT  14.0 3.2 14.8 14.8 ;
      RECT  2.8 6.6 3.6 7.4 ;
      RECT  7.6 8.6 8.4 9.4 ;
      RECT  1.2 5.2 2.0 10.8 ;
      RECT  18.8 9.4 19.6 10.2 ;
      RECT  7.6 8.6 8.4 9.4 ;
      RECT  35.8 6.1 36.4 6.7 ;
      RECT  30.2 12.1 30.8 12.7 ;
      RECT  2.8 6.6 3.6 7.4 ;
      RECT  4.4 36.8 5.2 25.2 ;
      RECT  14.0 36.8 14.8 25.2 ;
      RECT  2.8 33.4 3.6 32.6 ;
      RECT  7.6 31.4 8.4 30.6 ;
      RECT  1.2 34.8 2.0 29.2 ;
      RECT  18.8 30.6 19.6 29.8 ;
      RECT  7.6 31.4 8.4 30.6 ;
      RECT  35.8 33.9 36.4 33.3 ;
      RECT  30.2 27.9 30.8 27.3 ;
      RECT  2.8 33.4 3.6 32.6 ;
      RECT  7.6 8.6 8.4 9.4 ;
      RECT  7.6 30.6 8.4 31.4 ;
      RECT  35.8 6.1 36.4 6.7 ;
      RECT  30.2 12.1 30.8 12.7 ;
      RECT  35.8 33.3 36.4 33.9 ;
      RECT  30.2 27.3 30.8 27.9 ;
      RECT  2.8 0.0 3.4 40.0 ;
      RECT  31.4 162.8 30.8 172.4 ;
      RECT  3.1 162.8 2.5 329.2 ;
      RECT  7.6 8.6 8.4 9.4 ;
      RECT  7.6 30.6 8.4 31.4 ;
      RECT  51.7 9.5 52.3 10.1 ;
      RECT  30.8 162.8 31.4 172.4 ;
      RECT  63.5 150.1 77.0 150.7 ;
      RECT  63.3 88.7 77.0 89.3 ;
      RECT  69.1 109.9 77.0 110.5 ;
      RECT  70.9 70.7 77.0 71.3 ;
      RECT  72.4 8.7 77.0 9.3 ;
      RECT  59.6 345.2 60.4 356.8 ;
      RECT  69.2 345.2 70.0 356.8 ;
      RECT  58.0 348.6 58.8 349.4 ;
      RECT  62.8 350.6 63.6 351.4 ;
      RECT  56.4 347.2 57.2 352.8 ;
      RECT  74.0 351.4 74.8 352.2 ;
      RECT  59.6 378.8 60.4 367.2 ;
      RECT  69.2 378.8 70.0 367.2 ;
      RECT  58.0 375.4 58.8 374.6 ;
      RECT  62.8 373.4 63.6 372.6 ;
      RECT  56.4 376.8 57.2 371.2 ;
      RECT  74.0 372.6 74.8 371.8 ;
      RECT  59.6 385.2 60.4 396.8 ;
      RECT  69.2 385.2 70.0 396.8 ;
      RECT  58.0 388.6 58.8 389.4 ;
      RECT  62.8 390.6 63.6 391.4 ;
      RECT  56.4 387.2 57.2 392.8 ;
      RECT  74.0 391.4 74.8 392.2 ;
      RECT  59.6 418.8 60.4 407.2 ;
      RECT  69.2 418.8 70.0 407.2 ;
      RECT  58.0 415.4 58.8 414.6 ;
      RECT  62.8 413.4 63.6 412.6 ;
      RECT  56.4 416.8 57.2 411.2 ;
      RECT  74.0 412.6 74.8 411.8 ;
      RECT  62.8 350.6 63.6 351.4 ;
      RECT  62.8 372.6 63.6 373.4 ;
      RECT  62.8 390.6 63.6 391.4 ;
      RECT  62.8 412.6 63.6 413.4 ;
      RECT  74.0 351.4 74.8 352.2 ;
      RECT  74.0 371.8 74.8 372.6 ;
      RECT  74.0 391.4 74.8 392.2 ;
      RECT  74.0 411.8 74.8 412.6 ;
      RECT  103.2 34.2 104.0 45.8 ;
      RECT  112.8 34.2 113.6 45.8 ;
      RECT  101.6 37.6 102.4 38.4 ;
      RECT  106.4 39.6 107.2 40.4 ;
      RECT  100.0 36.2 100.8 41.8 ;
      RECT  117.6 40.4 118.4 41.2 ;
      RECT  125.0 34.2 125.8 45.8 ;
      RECT  134.6 34.2 135.4 45.8 ;
      RECT  123.4 37.6 124.2 38.4 ;
      RECT  128.2 39.6 129.0 40.4 ;
      RECT  121.8 36.2 122.6 41.8 ;
      RECT  139.4 40.4 140.2 41.2 ;
      RECT  106.4 39.6 107.2 40.4 ;
      RECT  128.2 39.6 129.0 40.4 ;
      RECT  117.6 40.4 118.4 41.2 ;
      RECT  139.4 40.4 140.2 41.2 ;
   LAYER  m3 ;
      RECT  180.7 172.8 181.5 173.6 ;
      RECT  180.7 360.0 181.5 360.8 ;
      RECT  177.3 167.8 178.1 168.6 ;
      RECT  184.1 355.0 184.9 355.8 ;
      RECT  184.1 167.8 184.9 168.6 ;
      RECT  177.3 355.0 178.1 355.8 ;
      RECT  173.9 256.0 174.7 256.8 ;
      RECT  173.9 235.2 174.7 236.0 ;
      RECT  201.1 256.0 201.9 256.8 ;
      RECT  173.9 318.4 174.7 319.2 ;
      RECT  180.7 360.0 181.5 360.8 ;
      RECT  201.1 172.8 201.9 173.6 ;
      RECT  201.1 193.6 201.9 194.4 ;
      RECT  201.1 360.0 201.9 360.8 ;
      RECT  173.9 360.0 174.7 360.8 ;
      RECT  173.9 193.6 174.7 194.4 ;
      RECT  173.9 297.6 174.7 298.4 ;
      RECT  201.1 214.4 201.9 215.2 ;
      RECT  173.9 214.4 174.7 215.2 ;
      RECT  187.5 360.0 188.3 360.8 ;
      RECT  194.3 360.0 195.1 360.8 ;
      RECT  180.7 172.8 181.5 173.6 ;
      RECT  201.1 318.4 201.9 319.2 ;
      RECT  173.9 339.2 174.7 340.0 ;
      RECT  187.5 172.8 188.3 173.6 ;
      RECT  173.9 172.8 174.7 173.6 ;
      RECT  201.1 235.2 201.9 236.0 ;
      RECT  194.3 172.8 195.1 173.6 ;
      RECT  201.1 339.2 201.9 340.0 ;
      RECT  201.1 297.6 201.9 298.4 ;
      RECT  201.1 276.8 201.9 277.6 ;
      RECT  173.9 276.8 174.7 277.6 ;
      RECT  184.1 167.8 184.9 168.6 ;
      RECT  184.1 167.8 184.9 168.6 ;
      RECT  177.3 313.4 178.1 314.2 ;
      RECT  177.3 271.8 178.1 272.6 ;
      RECT  204.5 355.0 205.3 355.8 ;
      RECT  170.5 240.2 171.3 241.0 ;
      RECT  170.5 302.6 171.3 303.4 ;
      RECT  204.5 344.2 205.3 345.0 ;
      RECT  177.3 177.8 178.1 178.6 ;
      RECT  197.7 188.6 198.5 189.4 ;
      RECT  177.3 198.6 178.1 199.4 ;
      RECT  170.5 313.4 171.3 314.2 ;
      RECT  170.5 271.8 171.3 272.6 ;
      RECT  170.5 167.8 171.3 168.6 ;
      RECT  204.5 292.6 205.3 293.4 ;
      RECT  177.3 219.4 178.1 220.2 ;
      RECT  197.7 219.4 198.5 220.2 ;
      RECT  197.7 334.2 198.5 335.0 ;
      RECT  204.5 334.2 205.3 335.0 ;
      RECT  170.5 344.2 171.3 345.0 ;
      RECT  170.5 355.0 171.3 355.8 ;
      RECT  197.7 292.6 198.5 293.4 ;
      RECT  197.7 355.0 198.5 355.8 ;
      RECT  197.7 177.8 198.5 178.6 ;
      RECT  170.5 323.4 171.3 324.2 ;
      RECT  197.7 271.8 198.5 272.6 ;
      RECT  170.5 219.4 171.3 220.2 ;
      RECT  204.5 177.8 205.3 178.6 ;
      RECT  204.5 281.8 205.3 282.6 ;
      RECT  177.3 292.6 178.1 293.4 ;
      RECT  197.7 344.2 198.5 345.0 ;
      RECT  170.5 251.0 171.3 251.8 ;
      RECT  204.5 302.6 205.3 303.4 ;
      RECT  204.5 240.2 205.3 241.0 ;
      RECT  170.5 230.2 171.3 231.0 ;
      RECT  204.5 188.6 205.3 189.4 ;
      RECT  197.7 261.0 198.5 261.8 ;
      RECT  177.3 251.0 178.1 251.8 ;
      RECT  197.7 167.8 198.5 168.6 ;
      RECT  177.3 334.2 178.1 335.0 ;
      RECT  197.7 323.4 198.5 324.2 ;
      RECT  170.5 292.6 171.3 293.4 ;
      RECT  197.7 251.0 198.5 251.8 ;
      RECT  177.3 167.8 178.1 168.6 ;
      RECT  177.3 167.8 178.1 168.6 ;
      RECT  204.5 209.4 205.3 210.2 ;
      RECT  170.5 188.6 171.3 189.4 ;
      RECT  177.3 209.4 178.1 210.2 ;
      RECT  204.5 198.6 205.3 199.4 ;
      RECT  177.3 344.2 178.1 345.0 ;
      RECT  170.5 334.2 171.3 335.0 ;
      RECT  197.7 302.6 198.5 303.4 ;
      RECT  177.3 281.8 178.1 282.6 ;
      RECT  204.5 261.0 205.3 261.8 ;
      RECT  197.7 313.4 198.5 314.2 ;
      RECT  190.9 167.8 191.7 168.6 ;
      RECT  170.5 261.0 171.3 261.8 ;
      RECT  204.5 230.2 205.3 231.0 ;
      RECT  190.9 355.0 191.7 355.8 ;
      RECT  177.3 188.6 178.1 189.4 ;
      RECT  197.7 281.8 198.5 282.6 ;
      RECT  204.5 271.8 205.3 272.6 ;
      RECT  184.1 355.0 184.9 355.8 ;
      RECT  170.5 209.4 171.3 210.2 ;
      RECT  184.1 355.0 184.9 355.8 ;
      RECT  170.5 177.8 171.3 178.6 ;
      RECT  177.3 230.2 178.1 231.0 ;
      RECT  177.3 240.2 178.1 241.0 ;
      RECT  197.7 209.4 198.5 210.2 ;
      RECT  197.7 230.2 198.5 231.0 ;
      RECT  197.7 198.6 198.5 199.4 ;
      RECT  170.5 198.6 171.3 199.4 ;
      RECT  197.7 240.2 198.5 241.0 ;
      RECT  204.5 167.8 205.3 168.6 ;
      RECT  204.5 323.4 205.3 324.2 ;
      RECT  204.5 313.4 205.3 314.2 ;
      RECT  177.3 302.6 178.1 303.4 ;
      RECT  204.5 251.0 205.3 251.8 ;
      RECT  177.3 355.0 178.1 355.8 ;
      RECT  177.3 355.0 178.1 355.8 ;
      RECT  170.5 281.8 171.3 282.6 ;
      RECT  177.3 323.4 178.1 324.2 ;
      RECT  177.3 261.0 178.1 261.8 ;
      RECT  204.5 219.4 205.3 220.2 ;
      RECT  181.2 156.8 182.0 157.6 ;
      RECT  188.0 156.8 188.8 157.6 ;
      RECT  194.8 156.8 195.6 157.6 ;
      RECT  181.2 156.8 182.0 157.6 ;
      RECT  188.0 156.8 188.8 157.6 ;
      RECT  194.8 156.8 195.6 157.6 ;
      RECT  189.9 122.6 190.7 123.4 ;
      RECT  196.7 122.6 197.5 123.4 ;
      RECT  197.7 136.0 198.5 136.8 ;
      RECT  190.9 136.0 191.7 136.8 ;
      RECT  195.1 71.2 195.9 72.0 ;
      RECT  194.5 88.6 195.3 89.4 ;
      RECT  187.7 88.6 188.5 89.4 ;
      RECT  188.3 71.2 189.1 72.0 ;
      RECT  189.7 82.2 190.5 83.0 ;
      RECT  195.1 77.8 195.9 78.6 ;
      RECT  196.5 82.2 197.3 83.0 ;
      RECT  193.7 96.8 194.5 97.6 ;
      RECT  188.3 77.8 189.1 78.6 ;
      RECT  186.9 96.8 187.7 97.6 ;
      RECT  189.9 123.4 190.7 122.6 ;
      RECT  188.3 72.0 189.1 71.2 ;
      RECT  181.2 157.6 182.0 156.8 ;
      RECT  196.7 123.4 197.5 122.6 ;
      RECT  187.7 89.4 188.5 88.6 ;
      RECT  194.8 157.6 195.6 156.8 ;
      RECT  188.0 157.6 188.8 156.8 ;
      RECT  194.5 89.4 195.3 88.6 ;
      RECT  195.1 72.0 195.9 71.2 ;
      RECT  188.3 78.6 189.1 77.8 ;
      RECT  196.5 83.0 197.3 82.2 ;
      RECT  193.7 97.6 194.5 96.8 ;
      RECT  197.7 136.8 198.5 136.0 ;
      RECT  195.1 78.6 195.9 77.8 ;
      RECT  186.9 97.6 187.7 96.8 ;
      RECT  190.9 136.8 191.7 136.0 ;
      RECT  189.7 83.0 190.5 82.2 ;
      RECT  90.7 214.8 91.5 215.6 ;
      RECT  105.7 214.8 106.5 215.6 ;
      RECT  105.7 214.8 106.5 215.6 ;
      RECT  90.7 194.0 91.5 194.8 ;
      RECT  105.7 194.0 106.5 194.8 ;
      RECT  105.7 194.0 106.5 194.8 ;
      RECT  90.7 194.0 91.5 194.8 ;
      RECT  90.7 214.8 91.5 215.6 ;
      RECT  105.7 183.6 106.5 184.4 ;
      RECT  90.7 225.2 91.5 226.0 ;
      RECT  105.7 204.4 106.5 205.2 ;
      RECT  90.7 183.6 91.5 184.4 ;
      RECT  90.7 204.4 91.5 205.2 ;
      RECT  105.7 225.2 106.5 226.0 ;
      RECT  90.7 277.2 91.5 278.0 ;
      RECT  105.7 277.2 106.5 278.0 ;
      RECT  105.7 277.2 106.5 278.0 ;
      RECT  90.7 256.4 91.5 257.2 ;
      RECT  105.7 256.4 106.5 257.2 ;
      RECT  105.7 256.4 106.5 257.2 ;
      RECT  90.7 256.4 91.5 257.2 ;
      RECT  90.7 277.2 91.5 278.0 ;
      RECT  105.7 246.0 106.5 246.8 ;
      RECT  90.7 287.6 91.5 288.4 ;
      RECT  105.7 266.8 106.5 267.6 ;
      RECT  90.7 246.0 91.5 246.8 ;
      RECT  90.7 266.8 91.5 267.6 ;
      RECT  105.7 287.6 106.5 288.4 ;
      RECT  90.7 194.0 91.5 194.8 ;
      RECT  90.7 277.2 91.5 278.0 ;
      RECT  149.6 277.2 150.4 278.0 ;
      RECT  149.6 256.4 150.4 257.2 ;
      RECT  149.6 214.8 150.4 215.6 ;
      RECT  149.6 214.8 150.4 215.6 ;
      RECT  149.6 256.4 150.4 257.2 ;
      RECT  149.6 194.0 150.4 194.8 ;
      RECT  105.7 256.4 106.5 257.2 ;
      RECT  90.7 214.8 91.5 215.6 ;
      RECT  105.7 277.2 106.5 278.0 ;
      RECT  105.7 214.8 106.5 215.6 ;
      RECT  90.7 256.4 91.5 257.2 ;
      RECT  149.6 194.0 150.4 194.8 ;
      RECT  149.6 235.6 150.4 236.4 ;
      RECT  149.6 298.0 150.4 298.8 ;
      RECT  149.6 318.8 150.4 319.6 ;
      RECT  149.6 339.6 150.4 340.4 ;
      RECT  149.6 277.2 150.4 278.0 ;
      RECT  105.7 194.0 106.5 194.8 ;
      RECT  90.7 183.6 91.5 184.4 ;
      RECT  105.7 266.8 106.5 267.6 ;
      RECT  90.7 246.0 91.5 246.8 ;
      RECT  149.6 350.0 150.4 350.8 ;
      RECT  90.7 204.4 91.5 205.2 ;
      RECT  105.7 287.6 106.5 288.4 ;
      RECT  90.7 225.2 91.5 226.0 ;
      RECT  105.7 204.4 106.5 205.2 ;
      RECT  105.7 225.2 106.5 226.0 ;
      RECT  149.6 246.0 150.4 246.8 ;
      RECT  149.6 287.6 150.4 288.4 ;
      RECT  105.7 183.6 106.5 184.4 ;
      RECT  90.7 287.6 91.5 288.4 ;
      RECT  149.6 225.2 150.4 226.0 ;
      RECT  149.6 204.4 150.4 205.2 ;
      RECT  105.7 246.0 106.5 246.8 ;
      RECT  149.6 266.8 150.4 267.6 ;
      RECT  149.6 329.2 150.4 330.0 ;
      RECT  149.6 308.4 150.4 309.2 ;
      RECT  149.6 183.6 150.4 184.4 ;
      RECT  90.7 266.8 91.5 267.6 ;
      RECT  165.1 235.6 165.9 236.4 ;
      RECT  165.1 298.0 165.9 298.8 ;
      RECT  165.1 256.4 165.9 257.2 ;
      RECT  165.1 256.4 165.9 257.2 ;
      RECT  165.1 277.2 165.9 278.0 ;
      RECT  165.1 277.2 165.9 278.0 ;
      RECT  165.1 214.8 165.9 215.6 ;
      RECT  165.1 214.8 165.9 215.6 ;
      RECT  165.1 194.0 165.9 194.8 ;
      RECT  165.1 194.0 165.9 194.8 ;
      RECT  165.1 339.6 165.9 340.4 ;
      RECT  165.1 318.8 165.9 319.6 ;
      RECT  165.1 350.0 165.9 350.8 ;
      RECT  165.1 246.0 165.9 246.8 ;
      RECT  165.1 225.2 165.9 226.0 ;
      RECT  165.1 329.2 165.9 330.0 ;
      RECT  165.1 183.6 165.9 184.4 ;
      RECT  165.1 266.8 165.9 267.6 ;
      RECT  165.1 204.4 165.9 205.2 ;
      RECT  165.1 287.6 165.9 288.4 ;
      RECT  165.1 308.4 165.9 309.2 ;
      RECT  165.1 318.8 165.9 319.6 ;
      RECT  90.7 256.4 91.5 257.2 ;
      RECT  165.1 298.0 165.9 298.8 ;
      RECT  165.1 277.2 165.9 278.0 ;
      RECT  149.6 235.6 150.4 236.4 ;
      RECT  149.6 214.8 150.4 215.6 ;
      RECT  105.7 277.2 106.5 278.0 ;
      RECT  149.6 298.0 150.4 298.8 ;
      RECT  90.7 214.8 91.5 215.6 ;
      RECT  105.7 194.0 106.5 194.8 ;
      RECT  165.1 194.0 165.9 194.8 ;
      RECT  165.1 339.6 165.9 340.4 ;
      RECT  165.1 214.8 165.9 215.6 ;
      RECT  149.6 339.6 150.4 340.4 ;
      RECT  165.1 256.4 165.9 257.2 ;
      RECT  149.6 194.0 150.4 194.8 ;
      RECT  90.7 194.0 91.5 194.8 ;
      RECT  105.7 214.8 106.5 215.6 ;
      RECT  149.6 256.4 150.4 257.2 ;
      RECT  149.6 318.8 150.4 319.6 ;
      RECT  105.7 256.4 106.5 257.2 ;
      RECT  90.7 277.2 91.5 278.0 ;
      RECT  165.1 235.6 165.9 236.4 ;
      RECT  149.6 277.2 150.4 278.0 ;
      RECT  105.7 266.8 106.5 267.6 ;
      RECT  105.7 204.4 106.5 205.2 ;
      RECT  149.6 183.6 150.4 184.4 ;
      RECT  90.7 246.0 91.5 246.8 ;
      RECT  149.6 266.8 150.4 267.6 ;
      RECT  105.7 183.6 106.5 184.4 ;
      RECT  149.6 350.0 150.4 350.8 ;
      RECT  165.1 225.2 165.9 226.0 ;
      RECT  105.7 287.6 106.5 288.4 ;
      RECT  90.7 287.6 91.5 288.4 ;
      RECT  90.7 266.8 91.5 267.6 ;
      RECT  165.1 183.6 165.9 184.4 ;
      RECT  90.7 183.6 91.5 184.4 ;
      RECT  105.7 246.0 106.5 246.8 ;
      RECT  165.1 308.4 165.9 309.2 ;
      RECT  165.1 329.2 165.9 330.0 ;
      RECT  165.1 204.4 165.9 205.2 ;
      RECT  149.6 308.4 150.4 309.2 ;
      RECT  149.6 246.0 150.4 246.8 ;
      RECT  149.6 225.2 150.4 226.0 ;
      RECT  165.1 287.6 165.9 288.4 ;
      RECT  165.1 350.0 165.9 350.8 ;
      RECT  90.7 204.4 91.5 205.2 ;
      RECT  149.6 204.4 150.4 205.2 ;
      RECT  165.1 266.8 165.9 267.6 ;
      RECT  149.6 329.2 150.4 330.0 ;
      RECT  90.7 225.2 91.5 226.0 ;
      RECT  165.1 246.0 165.9 246.8 ;
      RECT  149.6 287.6 150.4 288.4 ;
      RECT  105.7 225.2 106.5 226.0 ;
      RECT  173.9 256.0 174.7 256.8 ;
      RECT  165.1 277.2 165.9 278.0 ;
      RECT  195.1 71.2 195.9 72.0 ;
      RECT  165.1 339.6 165.9 340.4 ;
      RECT  173.9 235.2 174.7 236.0 ;
      RECT  201.1 256.0 201.9 256.8 ;
      RECT  181.2 156.8 182.0 157.6 ;
      RECT  90.7 214.8 91.5 215.6 ;
      RECT  173.9 318.4 174.7 319.2 ;
      RECT  180.7 360.0 181.5 360.8 ;
      RECT  201.1 172.8 201.9 173.6 ;
      RECT  201.1 193.6 201.9 194.4 ;
      RECT  149.6 277.2 150.4 278.0 ;
      RECT  201.1 360.0 201.9 360.8 ;
      RECT  173.9 360.0 174.7 360.8 ;
      RECT  173.9 193.6 174.7 194.4 ;
      RECT  173.9 297.6 174.7 298.4 ;
      RECT  201.1 214.4 201.9 215.2 ;
      RECT  173.9 214.4 174.7 215.2 ;
      RECT  189.9 122.6 190.7 123.4 ;
      RECT  149.6 194.0 150.4 194.8 ;
      RECT  90.7 194.0 91.5 194.8 ;
      RECT  105.7 214.8 106.5 215.6 ;
      RECT  149.6 298.0 150.4 298.8 ;
      RECT  149.6 256.4 150.4 257.2 ;
      RECT  194.5 88.6 195.3 89.4 ;
      RECT  187.5 360.0 188.3 360.8 ;
      RECT  194.3 360.0 195.1 360.8 ;
      RECT  180.7 172.8 181.5 173.6 ;
      RECT  201.1 318.4 201.9 319.2 ;
      RECT  196.7 122.6 197.5 123.4 ;
      RECT  188.3 71.2 189.1 72.0 ;
      RECT  105.7 277.2 106.5 278.0 ;
      RECT  165.1 214.8 165.9 215.6 ;
      RECT  165.1 298.0 165.9 298.8 ;
      RECT  194.8 156.8 195.6 157.6 ;
      RECT  187.7 88.6 188.5 89.4 ;
      RECT  165.1 194.0 165.9 194.8 ;
      RECT  90.7 277.2 91.5 278.0 ;
      RECT  90.7 256.4 91.5 257.2 ;
      RECT  149.6 214.8 150.4 215.6 ;
      RECT  173.9 339.2 174.7 340.0 ;
      RECT  165.1 256.4 165.9 257.2 ;
      RECT  187.5 172.8 188.3 173.6 ;
      RECT  188.0 156.8 188.8 157.6 ;
      RECT  149.6 235.6 150.4 236.4 ;
      RECT  173.9 172.8 174.7 173.6 ;
      RECT  165.1 318.8 165.9 319.6 ;
      RECT  165.1 235.6 165.9 236.4 ;
      RECT  201.1 235.2 201.9 236.0 ;
      RECT  105.7 256.4 106.5 257.2 ;
      RECT  194.3 172.8 195.1 173.6 ;
      RECT  149.6 318.8 150.4 319.6 ;
      RECT  201.1 339.2 201.9 340.0 ;
      RECT  201.1 297.6 201.9 298.4 ;
      RECT  149.6 339.6 150.4 340.4 ;
      RECT  105.7 194.0 106.5 194.8 ;
      RECT  201.1 276.8 201.9 277.6 ;
      RECT  173.9 276.8 174.7 277.6 ;
      RECT  184.1 167.8 184.9 168.6 ;
      RECT  177.3 313.4 178.1 314.2 ;
      RECT  90.7 266.8 91.5 267.6 ;
      RECT  177.3 271.8 178.1 272.6 ;
      RECT  204.5 355.0 205.3 355.8 ;
      RECT  170.5 240.2 171.3 241.0 ;
      RECT  170.5 302.6 171.3 303.4 ;
      RECT  204.5 344.2 205.3 345.0 ;
      RECT  177.3 177.8 178.1 178.6 ;
      RECT  197.7 188.6 198.5 189.4 ;
      RECT  177.3 198.6 178.1 199.4 ;
      RECT  170.5 313.4 171.3 314.2 ;
      RECT  165.1 204.4 165.9 205.2 ;
      RECT  170.5 271.8 171.3 272.6 ;
      RECT  188.3 77.8 189.1 78.6 ;
      RECT  149.6 246.0 150.4 246.8 ;
      RECT  170.5 167.8 171.3 168.6 ;
      RECT  204.5 292.6 205.3 293.4 ;
      RECT  177.3 219.4 178.1 220.2 ;
      RECT  149.6 225.2 150.4 226.0 ;
      RECT  165.1 246.0 165.9 246.8 ;
      RECT  197.7 219.4 198.5 220.2 ;
      RECT  105.7 183.6 106.5 184.4 ;
      RECT  197.7 334.2 198.5 335.0 ;
      RECT  204.5 334.2 205.3 335.0 ;
      RECT  149.6 266.8 150.4 267.6 ;
      RECT  149.6 204.4 150.4 205.2 ;
      RECT  170.5 344.2 171.3 345.0 ;
      RECT  170.5 355.0 171.3 355.8 ;
      RECT  197.7 292.6 198.5 293.4 ;
      RECT  197.7 355.0 198.5 355.8 ;
      RECT  197.7 177.8 198.5 178.6 ;
      RECT  170.5 323.4 171.3 324.2 ;
      RECT  197.7 271.8 198.5 272.6 ;
      RECT  170.5 219.4 171.3 220.2 ;
      RECT  204.5 177.8 205.3 178.6 ;
      RECT  204.5 281.8 205.3 282.6 ;
      RECT  90.7 287.6 91.5 288.4 ;
      RECT  177.3 292.6 178.1 293.4 ;
      RECT  186.9 96.8 187.7 97.6 ;
      RECT  165.1 350.0 165.9 350.8 ;
      RECT  197.7 344.2 198.5 345.0 ;
      RECT  170.5 251.0 171.3 251.8 ;
      RECT  204.5 302.6 205.3 303.4 ;
      RECT  105.7 287.6 106.5 288.4 ;
      RECT  204.5 240.2 205.3 241.0 ;
      RECT  170.5 230.2 171.3 231.0 ;
      RECT  149.6 183.6 150.4 184.4 ;
      RECT  165.1 266.8 165.9 267.6 ;
      RECT  204.5 188.6 205.3 189.4 ;
      RECT  197.7 261.0 198.5 261.8 ;
      RECT  177.3 251.0 178.1 251.8 ;
      RECT  197.7 167.8 198.5 168.6 ;
      RECT  193.7 96.8 194.5 97.6 ;
      RECT  177.3 334.2 178.1 335.0 ;
      RECT  197.7 323.4 198.5 324.2 ;
      RECT  170.5 292.6 171.3 293.4 ;
      RECT  197.7 251.0 198.5 251.8 ;
      RECT  177.3 167.8 178.1 168.6 ;
      RECT  204.5 209.4 205.3 210.2 ;
      RECT  170.5 188.6 171.3 189.4 ;
      RECT  177.3 209.4 178.1 210.2 ;
      RECT  204.5 198.6 205.3 199.4 ;
      RECT  149.6 329.2 150.4 330.0 ;
      RECT  197.7 136.0 198.5 136.8 ;
      RECT  195.1 77.8 195.9 78.6 ;
      RECT  177.3 344.2 178.1 345.0 ;
      RECT  170.5 334.2 171.3 335.0 ;
      RECT  105.7 266.8 106.5 267.6 ;
      RECT  90.7 183.6 91.5 184.4 ;
      RECT  197.7 302.6 198.5 303.4 ;
      RECT  177.3 281.8 178.1 282.6 ;
      RECT  204.5 261.0 205.3 261.8 ;
      RECT  197.7 313.4 198.5 314.2 ;
      RECT  165.1 329.2 165.9 330.0 ;
      RECT  190.9 167.8 191.7 168.6 ;
      RECT  105.7 225.2 106.5 226.0 ;
      RECT  165.1 308.4 165.9 309.2 ;
      RECT  170.5 261.0 171.3 261.8 ;
      RECT  204.5 230.2 205.3 231.0 ;
      RECT  165.1 287.6 165.9 288.4 ;
      RECT  190.9 355.0 191.7 355.8 ;
      RECT  177.3 188.6 178.1 189.4 ;
      RECT  197.7 281.8 198.5 282.6 ;
      RECT  149.6 308.4 150.4 309.2 ;
      RECT  204.5 271.8 205.3 272.6 ;
      RECT  90.7 225.2 91.5 226.0 ;
      RECT  184.1 355.0 184.9 355.8 ;
      RECT  170.5 209.4 171.3 210.2 ;
      RECT  90.7 246.0 91.5 246.8 ;
      RECT  149.6 350.0 150.4 350.8 ;
      RECT  170.5 177.8 171.3 178.6 ;
      RECT  177.3 230.2 178.1 231.0 ;
      RECT  105.7 204.4 106.5 205.2 ;
      RECT  165.1 225.2 165.9 226.0 ;
      RECT  177.3 240.2 178.1 241.0 ;
      RECT  197.7 209.4 198.5 210.2 ;
      RECT  197.7 230.2 198.5 231.0 ;
      RECT  197.7 198.6 198.5 199.4 ;
      RECT  170.5 198.6 171.3 199.4 ;
      RECT  197.7 240.2 198.5 241.0 ;
      RECT  190.9 136.0 191.7 136.8 ;
      RECT  204.5 167.8 205.3 168.6 ;
      RECT  149.6 287.6 150.4 288.4 ;
      RECT  204.5 323.4 205.3 324.2 ;
      RECT  90.7 204.4 91.5 205.2 ;
      RECT  204.5 313.4 205.3 314.2 ;
      RECT  177.3 302.6 178.1 303.4 ;
      RECT  204.5 251.0 205.3 251.8 ;
      RECT  177.3 355.0 178.1 355.8 ;
      RECT  105.7 246.0 106.5 246.8 ;
      RECT  170.5 281.8 171.3 282.6 ;
      RECT  196.5 82.2 197.3 83.0 ;
      RECT  189.7 82.2 190.5 83.0 ;
      RECT  177.3 323.4 178.1 324.2 ;
      RECT  177.3 261.0 178.1 261.8 ;
      RECT  204.5 219.4 205.3 220.2 ;
      RECT  165.1 183.6 165.9 184.4 ;
      RECT  -0.4 19.6 0.4 20.4 ;
      RECT  -0.4 39.6 0.4 40.4 ;
      RECT  -0.4 -0.4 0.4 0.4 ;
      RECT  8.4 182.0 7.6 182.8 ;
      RECT  21.6 221.2 20.8 222.0 ;
      RECT  8.4 260.4 7.6 261.2 ;
      RECT  8.4 221.2 7.6 222.0 ;
      RECT  8.4 299.6 7.6 300.4 ;
      RECT  21.6 299.6 20.8 300.4 ;
      RECT  8.4 338.8 7.6 339.6 ;
      RECT  21.6 182.0 20.8 182.8 ;
      RECT  21.6 260.4 20.8 261.2 ;
      RECT  21.6 338.8 20.8 339.6 ;
      RECT  21.6 319.2 20.8 320.0 ;
      RECT  8.4 201.6 7.6 202.4 ;
      RECT  8.4 280.0 7.6 280.8 ;
      RECT  21.6 280.0 20.8 280.8 ;
      RECT  8.4 162.4 7.6 163.2 ;
      RECT  21.6 240.8 20.8 241.6 ;
      RECT  8.4 319.2 7.6 320.0 ;
      RECT  21.6 162.4 20.8 163.2 ;
      RECT  8.4 240.8 7.6 241.6 ;
      RECT  21.6 201.6 20.8 202.4 ;
      RECT  20.8 260.4 21.6 261.2 ;
      RECT  7.6 338.8 8.4 339.6 ;
      RECT  7.6 182.0 8.4 182.8 ;
      RECT  75.2 19.6 76.0 20.4 ;
      RECT  7.6 221.2 8.4 222.0 ;
      RECT  75.2 139.6 76.0 140.4 ;
      RECT  75.2 59.6 76.0 60.4 ;
      RECT  20.8 182.0 21.6 182.8 ;
      RECT  7.6 260.4 8.4 261.2 ;
      RECT  7.6 299.6 8.4 300.4 ;
      RECT  -0.4 19.6 0.4 20.4 ;
      RECT  20.8 338.8 21.6 339.6 ;
      RECT  20.8 221.2 21.6 222.0 ;
      RECT  20.8 299.6 21.6 300.4 ;
      RECT  75.2 99.6 76.0 100.4 ;
      RECT  75.2 119.6 76.0 120.4 ;
      RECT  20.8 280.0 21.6 280.8 ;
      RECT  -0.4 -0.4 0.4 0.4 ;
      RECT  75.2 159.6 76.0 160.4 ;
      RECT  20.8 319.2 21.6 320.0 ;
      RECT  7.6 319.2 8.4 320.0 ;
      RECT  20.8 201.6 21.6 202.4 ;
      RECT  -0.4 39.6 0.4 40.4 ;
      RECT  75.2 39.6 76.0 40.4 ;
      RECT  7.6 201.6 8.4 202.4 ;
      RECT  75.2 -0.4 76.0 0.4 ;
      RECT  20.8 240.8 21.6 241.6 ;
      RECT  75.2 79.6 76.0 80.4 ;
      RECT  7.6 240.8 8.4 241.6 ;
      RECT  7.6 280.0 8.4 280.8 ;
      RECT  7.6 162.4 8.4 163.2 ;
      RECT  20.8 162.4 21.6 163.2 ;
      RECT  55.2 345.1 77.0 345.7 ;
      RECT  65.7 401.6 66.5 402.4 ;
      RECT  65.7 361.6 66.5 362.4 ;
      RECT  65.7 421.6 66.5 422.4 ;
      RECT  65.7 341.6 66.5 342.4 ;
      RECT  65.7 381.6 66.5 382.4 ;
      RECT  98.8 34.1 142.4 34.7 ;
      RECT  131.1 50.6 131.9 51.4 ;
      RECT  109.3 50.6 110.1 51.4 ;
      RECT  131.1 30.6 131.9 31.4 ;
      RECT  109.3 30.6 110.1 31.4 ;
   LAYER  m4 ;
   END
   END    sram_2_16_scn4m_subm
END    LIBRARY
